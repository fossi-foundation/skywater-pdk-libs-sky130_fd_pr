* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

******************************************************************
******************************************************************
*  *****************************************************
*  04/26/2021 Usman Suriono
*      Why     : New scalable sky130_fd_pr__nfet_01v8 VHV model
*      What    : Converted from discrete nvhv models
*                Changed the parasitic diode from internal dimension calculation
*                to receive it from PDK
*
*  *****************************************************
*
*  Nmos VHV DE Model
*  -----------------------------------------------------

.subckt  sky130_fd_pr__nfet_g5v0d16v0 d g s b mult=1
+ 
.param  w = 5 l = 0.7 nf = 1 sa = 0 sb = 0 sd = 0
*** All values are estimated, the real values supplied and overwritten by PDK netlist
+ ad = {3.89*(w+1.3)}
+ pd = {2*(3.89+w+1.3)}
+ as = {0.28*w}
+ ps = {2*(0.28+w)}
+ nrd = {0.135*nf/w}
+ nrs = {0.140*nf/w}


rldd d d1  r = {(1/w)*5906.5*sw_nw_rs_mult*1.03} tc1 = 1.483e-3 tc2 = 7.824e-6
xdnw1 b d sky130_fd_pr__model__parasitic__diode_pd2nw area = {ad} perim = {pd} m = 0.5
xdnw2 b d1 sky130_fd_pr__model__parasitic__diode_pd2nw area = {ad} perim = {pd} m = 0.5
Xsky130_fd_pr__nfet_g5v0d16v0 d1 g s b sky130_fd_pr__nfet_g5v0d16v0_base l = {l} w = {w} ad = 0 as = {as} pd = 0 ps = {ps} nrd = {nrd} nrs = {nrs*sw_rdn/sw_rnw} sa = {sa} sb = {sb} sd = {sd} nf = {nf}



.ends sky130_fd_pr__nfet_g5v0d16v0
