* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

*  -----------------------------------------------------
*       Base Nmos VHV DE Model
*  -----------------------------------------------------

.subckt  sky130_fd_pr__nfet_g5v0d16v0_base  d g s b  mult=1
+ l=1 w=1 
.param  nf = 1 ad = 0 as = 0 pd = 0 ps = 0 nrd = 0 nrs = 0 sa = 0 sb = 0 sd = 0
+ swx_vth0_delta = {sw_vth0_sky130_fd_pr__nfet_g5v0d16v0+sw_mm_vth0_sky130_fd_pr__nfet_g5v0d16v0*mismatch_factor*MC_MM_SWITCH*AGAUSS(0,1.0,1)/sqrt(l*w*mult)+sw_vth0_sky130_fd_pr__nfet_g5v0d16v0_mc}


Msky130_fd_pr__nfet_g5v0d16v0_base  d g s b nvhv_model_base l = {l} w = {w} ad = {ad} as = {as} pd = {pd} ps = {ps} nrd = {nrd} nrs = {nrs} sa = {sa} sb = {sb} sd = {sd} nf = {nf}
* + deltox = 0.3*(sw_tox_hv_corner - sw_tox_hv_nom) + sw_tox_hv_mc + sw_mm_tox_hv * mismatch_factor*MC_MM_SWITCH*AGAUSS(0,1.0,1)/sqrt(l*w*mult)
* + mulu0  = sw_u0_sky130_fd_pr__nfet_g5v0d16v0
+ delvto = {-0.0005+swx_vth0_delta*(0.090*2.2/l+0.91)*(0.0005*44/(w*l)+0.9995)}
* + delk1  = 0.27 * swx_vth0_delta
* + mulvsat = sw_vsat_sky130_fd_pr__nfet_g5v0d16v0




.model nvhv_model_base.1 nmos
+ level = 54 lmin = 2.2E-6 lmax = 2.02E-5 wmin = 6E-5
+ wmax = 1.01E-3 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 1 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 1.16E-8
+ toxm = 1.16E-8 xj = 1.5E-7 ndep = 1.7E17
+ ngate = 1E23 nsd = 1E20 rsh = {sw_rnw}
+ rshg = 0.1 phin = 0 wint = {2.1346E-8+sw_activecd}
+ wl = 0 wln = 1 ww = 0
+ wwn = 1 wwl = 0 lint = {7.6507E-8-sw_polycd}
+ ll = 0 lln = 1 lw = 0
+ lwn = 1 lwl = 0 llc = 0
+ lwc = 0 lwlc = 0 wlc = 0
+ wwc = 0 wwlc = 0 dwg = -4.1292E-9
+ dwb = -1.6944E-9 xl = 0 xw = 0
+ dmcg = 0 dmdg = 0 dmcgt = 0
+ xgw = 0 xgl = 0 ngcon = 1
+ vth0 = 0.795183 k1 = 0.89738 k2 = -0.044197
+ k3 = -0.884 k3b = 0.43 w0 = 0
+ lpe0 = 0 lpeb = -2.182E-7 vbm = -3
+ dvtp0 = 0 dvtp1 = 0 dvt0 = 0
+ dvt1 = 0.53 dvt2 = -0.19251 dvt0w = 0.16
+ dvt1w = 6.9091E6 dvt2w = -0.036016 u0 = 3.54241E-2
+ ua = 8E-11 ub = 2.1405E-18 uc = 6.0747E-11
+ ud = 0 up = 0 lp = 1
+ eu = 1.67 vsat = 1.0055E5 a0 = 0.3
+ ags = 0.13326 b0 = 3.2933E-8 b1 = 0
+ keta = -0.05 a1 = 0 a2 = 0.659726
+ rdsw = 724.62 rdswmin = 0 rdw = 1
+ rdwmin = 0 rsw = 0 rswmin = 0
+ prwb = 0 prwg = 0 wr = 1
+ voff = -0.20613 voffl = -4.257949E-7 minv = 0
+ nfactor = 0.83837 eta0 = 0.016128 etab = -0.02983
+ dsub = 0.504 cit = -8E-4 cdsc = 0
+ cdscb = 0 cdscd = 0 pclm = 0.16548
+ pdiblc1 = 0.21098 pdiblc2 = 2E-4 pdiblcb = -0.26831
+ drout = 0.36652 pscbe1 = 9.3731E8 pscbe2 = 1.68E-6
+ pvag = 1.99 delta = 1E-3 fprout = 10.125
+ pdits = 0 pditsl = 0 pditsd = 0
+ vtl = 0 xn = 3 alpha0 = 3.0448E-7
+ alpha1 = 0.72 beta0 = 37.72 aigbacc = 1
+ bigbacc = 0 cigbacc = 0 nigbacc = 1
+ aigbinv = 0.35 bigbinv = 0.03 cigbinv = 6E-3
+ eigbinv = 1.1 nigbinv = 3 aigc = 0.43
+ bigc = 0.054 cigc = 0.075 aigsd = 0.43
+ bigsd = 0.054 cigsd = 0.075 dlcig = 0
+ nigc = 1 poxedge = 1 pigcd = 1
+ ntox = 1 toxref = 1.16E-8 agidl = 0
+ bgidl = 1.058E9 cgidl = 4E3 egidl = 0.8
+ noia = 2.6E41 noib = 0 noic = 0
+ em = 4.1E7 ef = 0.89 lintnoi = 0
+ tnoia = 7.5E6 tnoib = 7.2E6 rnoia = 0.794
+ rnoib = 0.38 xpart = 0 cgso = {1.5674E-10/sw_func_tox_hv_ratio}
+ cgdo = {3.0674E-10/sw_func_tox_hv_ratio} cgbo = {0/sw_func_tox_hv_ratio} ckappas = 0.6
+ cf = 0 clc = 1E-7 cle = 0.6
+ dlc = -3.5995E-8 dwc = 0 vfbcv = -1
+ noff = 4 voffcv = -0.2104 acde = 0.4176
+ moin = 15 cgsl = {4.49025E-11/sw_func_tox_hv_ratio} cgdl = {4.49025E-11/sw_func_tox_hv_ratio}
+ ijthsrev = 0.1 ijthsfwd = 0.1 xjbvs = 1
+ bvs = 12.636 jss = 3.75E-4 jsws = 5.84E-11
+ cjs = {8.310E-04*sw_func_nsd_pw_cj} mjs = 0.295 mjsws = 0.037586
+ cjsws = {8.643094E-11*sw_func_nsd_pw_cj} cjswgs = {5.47776E-11*sw_func_nsd_pw_cj} mjswgs = 0.78692
+ pbs = 0.72468 pbsws = 0.29067 pbswgs = 0.54958
+ tnom = 30 ute = -1.4324 kt1 = -0.37073
+ kt1l = 0 kt2 = -0.019151 ua1 = 2.0117E-9
+ ub1 = -2.9862E-18 uc1 = -5.9821E-11 at = 2.9E4
+ prt = 0 njs = 1.0773 xtis = 0.76
+ tpb = 1.344E-3 tpbsw = 9.9005E-4 tpbswg = 0
+ tcj = 6.7434E-4 tcjsw = 2.493E-4 tcjswg = 0
+ tvoff = 0 saref = 2.8E-7 sbref = 1.585E-6
+ wlod = 0 ku0 = -9.9E-8 kvsat = 0.3
+ kvth0 = 1.7057E-8 tku0 = 0 llodku0 = 1
+ wlodku0 = 1 llodvth = 1 wlodvth = 1
+ lku0 = 9.6975E-7 wku0 = 2E-7 pku0 = 0
+ lkvth0 = 2.2691E-7 wkvth0 = 2.3093E-6 pkvth0 = 0
+ stk2 = 0 lodk2 = 1 steta0 = 0
+ lodeta0 = 1

.model nvhv_model_base.2 nmos
+ level = 54 lmin = 7E-7 lmax = 2.2E-6 wmin = 6E-5
+ wmax = 1.01E-3 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 1 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 1.16E-8
+ toxm = 1.16E-8 xj = 1.5E-7 ndep = 1.7E17
+ ngate = 1E23 nsd = 1E20 rsh = {sw_rnw}
+ rshg = 0.1 phin = 0 wint = {2.1346E-8+sw_activecd}
+ wl = 0 wln = 1 ww = 0
+ wwn = 1 wwl = 0 lint = {7.6507E-8-sw_polycd}
+ ll = 0 lln = 1 lw = 0
+ lwn = 1 lwl = 0 llc = 0
+ lwc = 0 lwlc = 0 wlc = 0
+ wwc = 0 wwlc = 0 dwg = -4.1292E-9
+ dwb = -1.6944E-9 xl = 0 xw = 0
+ dmcg = 0 dmdg = 0 dmcgt = 0
+ xgw = 0 xgl = 0 ngcon = 1
+ vth0 = 0.800438 lvth0 = -1.075632E-8 k1 = 0.923559
+ lk1 = -5.358753E-8 k2 = -4.92657E-2 lk2 = 1.037563E-8
+ k3 = -0.884 k3b = 0.43 w0 = 0
+ lpe0 = 0 lpeb = -2.182E-7 vbm = -3
+ dvtp0 = 0 dvtp1 = 0 dvt0 = 0
+ dvt1 = 0.53 dvt2 = -0.19251 dvt0w = 0.16
+ dvt1w = 6.9091E6 dvt2w = -0.036016 u0 = 3.39297E-2
+ lu0 = 3.059095E-9 ua = -9.595287E-10 lua = 2.127901E-15
+ ub = 2.645044E-18 lub = -1.032794E-24 uc = 7.074156E-11
+ luc = -2.045873E-17 ud = 0 up = 0
+ lp = 1 eu = 1.67 vsat = 1.104359E5
+ lvsat = -2.02362E-2 a0 = 0.141473 la0 = 3.245035E-7
+ ags = -0.198265 lags = 6.786261E-7 b0 = 3.2933E-8
+ b1 = 0 keta = 1.43127E-3 lketa = -1.052791E-7
+ a1 = 0 a2 = 0.659726 rdsw = 724.62
+ rdswmin = 0 rdw = 1 rdwmin = 0
+ rsw = 0 rswmin = 0 prwb = 0
+ prwg = 0 wr = 1 voff = -0.20613
+ voffl = -4.257949E-7 minv = 0 nfactor = 0.83837
+ eta0 = 0.016128 etab = -0.02983 dsub = 0.504
+ cit = -8E-4 cdsc = 0 cdscb = 0
+ cdscd = 0 pclm = -7.58976E-2 lpclm = 4.940966E-7
+ pdiblc1 = 0.21098 pdiblc2 = 2E-4 pdiblcb = -0.26831
+ drout = 0.36652 pscbe1 = 9.3731E8 pscbe2 = 1.68E-6
+ pvag = 1.99 delta = -4.586293E-4 ldelta = 2.985794E-9
+ fprout = 10.125 pdits = 0 pditsl = 0
+ pditsd = 0 vtl = 0 xn = 3
+ alpha0 = -1.062595E-5 lalpha0 = 2.237443E-11 alpha1 = 0.573481
+ lalpha1 = 2.99923E-7 beta0 = 24.125575 lbeta0 = 2.78276E-5
+ aigbacc = 1 bigbacc = 0 cigbacc = 0
+ nigbacc = 1 aigbinv = 0.35 bigbinv = 0.03
+ cigbinv = 6E-3 eigbinv = 1.1 nigbinv = 3
+ aigc = 0.43 bigc = 0.054 cigc = 0.075
+ aigsd = 0.43 bigsd = 0.054 cigsd = 0.075
+ dlcig = 0 nigc = 1 poxedge = 1
+ pigcd = 1 ntox = 1 toxref = 1.16E-8
+ agidl = 0 bgidl = 1.058E9 cgidl = 4E3
+ egidl = 0.8 noia = 2.6E41 noib = 0
+ noic = 0 em = 4.1E7 ef = 0.89
+ lintnoi = 0 tnoia = 7.5E6 tnoib = 7.2E6
+ rnoia = 0.794 rnoib = 0.38 xpart = 0
+ cgso = {1.5674E-10/sw_func_tox_hv_ratio} cgdo = {3.0674E-10/sw_func_tox_hv_ratio} cgbo = {0/sw_func_tox_hv_ratio}
+ ckappas = 0.6 cf = 0 clc = 1E-7
+ cle = 0.6 dlc = -3.5995E-8 dwc = 0
+ vfbcv = -1 noff = 4 voffcv = -0.2104
+ acde = 0.4176 moin = 15 cgsl = {4.49025E-11/sw_func_tox_hv_ratio}
+ cgdl = {4.49025E-11/sw_func_tox_hv_ratio} ijthsrev = 0.1 ijthsfwd = 0.1
+ xjbvs = 1 bvs = 12.636 jss = 3.75E-4
+ jsws = 5.84E-11 cjs = {8.310E-04*sw_func_nsd_pw_cj} mjs = 0.295
+ mjsws = 0.037586 cjsws = {8.643094E-11*sw_func_nsd_pw_cj} cjswgs = {5.47776E-11*sw_func_nsd_pw_cj}
+ mjswgs = 0.78692 pbs = 0.72468 pbsws = 0.29067
+ pbswgs = 0.54958 tnom = 30 ute = -1.417741
+ lute = -3.000723E-8 kt1 = -0.37073 kt1l = 0
+ kt2 = -3.181197E-3 lkt2 = -3.268996E-8 ua1 = 2.0117E-9
+ ub1 = -3.237121E-18 lub1 = 5.136312E-25 uc1 = -8.080006E-11
+ luc1 = 4.294385E-17 at = 2.9E4 prt = 0
+ njs = 1.0773 xtis = 0.76 tpb = 1.344E-3
+ tpbsw = 9.9005E-4 tpbswg = 0 tcj = 6.7434E-4
+ tcjsw = 2.493E-4 tcjswg = 0 tvoff = 0
+ saref = 2.8E-7 sbref = 1.585E-6 wlod = 0
+ ku0 = -9.9E-8 kvsat = 0.3 kvth0 = 1.7057E-8
+ tku0 = 0 llodku0 = 1 wlodku0 = 1
+ llodvth = 1 wlodvth = 1 lku0 = 9.6975E-7
+ wku0 = 2E-7 pku0 = 0 lkvth0 = 2.2691E-7
+ wkvth0 = 2.3093E-6 pkvth0 = 0 stk2 = 0
+ lodk2 = 1 steta0 = 0 lodeta0 = 1

.model nvhv_model_base.3 nmos
+ level = 54 lmin = 2.2E-6 lmax = 2.02E-5 wmin = 5E-5
+ wmax = 6E-5 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 1 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 1.16E-8
+ toxm = 1.16E-8 xj = 1.5E-7 ndep = 1.7E17
+ ngate = 1E23 nsd = 1E20 rsh = {sw_rnw}
+ rshg = 0.1 phin = 0 wint = {2.1346E-8+sw_activecd}
+ wl = 0 wln = 1 ww = 0
+ wwn = 1 wwl = 0 lint = {7.6507E-8-sw_polycd}
+ ll = 0 lln = 1 lw = 0
+ lwn = 1 lwl = 0 llc = 0
+ lwc = 0 lwlc = 0 wlc = 0
+ wwc = 0 wwlc = 0 dwg = -4.1292E-9
+ dwb = -1.6944E-9 xl = 0 xw = 0
+ dmcg = 0 dmdg = 0 dmcgt = 0
+ xgw = 0 xgl = 0 ngcon = 1
+ vth0 = 0.795183 k1 = 0.89738 k2 = -0.044197
+ k3 = -0.884 k3b = 0.43 w0 = 0
+ lpe0 = 0 lpeb = -2.182E-7 vbm = -3
+ dvtp0 = 0 dvtp1 = 0 dvt0 = 0
+ dvt1 = 0.53 dvt2 = -0.19251 dvt0w = 0.16
+ dvt1w = 6.9091E6 dvt2w = -0.036016 u0 = 3.54241E-2
+ ua = 8E-11 ub = 2.1405E-18 uc = 6.0747E-11
+ ud = 0 up = 0 lp = 1
+ eu = 1.67 vsat = 1.0055E5 a0 = 0.3
+ ags = 0.13326 b0 = 3.2933E-8 b1 = 0
+ keta = -0.05 a1 = 0 a2 = 0.659726
+ rdsw = 724.62 rdswmin = 0 rdw = 1
+ rdwmin = 0 rsw = 0 rswmin = 0
+ prwb = 0 prwg = 0 wr = 1
+ voff = -0.20613 voffl = -4.257949E-7 minv = 0
+ nfactor = 0.83837 eta0 = 0.016128 etab = -0.02983
+ dsub = 0.504 cit = -8E-4 cdsc = 0
+ cdscb = 0 cdscd = 0 pclm = 0.16548
+ pdiblc1 = 0.21098 pdiblc2 = 2E-4 pdiblcb = -0.26831
+ drout = 0.36652 pscbe1 = 9.3731E8 pscbe2 = 1.68E-6
+ pvag = 1.99 delta = 1E-3 fprout = 10.125
+ pdits = 0 pditsl = 0 pditsd = 0
+ vtl = 0 xn = 3 alpha0 = 3.0448E-7
+ alpha1 = 0.72 beta0 = 37.72 aigbacc = 1
+ bigbacc = 0 cigbacc = 0 nigbacc = 1
+ aigbinv = 0.35 bigbinv = 0.03 cigbinv = 6E-3
+ eigbinv = 1.1 nigbinv = 3 aigc = 0.43
+ bigc = 0.054 cigc = 0.075 aigsd = 0.43
+ bigsd = 0.054 cigsd = 0.075 dlcig = 0
+ nigc = 1 poxedge = 1 pigcd = 1
+ ntox = 1 toxref = 1.16E-8 agidl = 0
+ bgidl = 1.058E9 cgidl = 4E3 egidl = 0.8
+ noia = 2.6E41 noib = 0 noic = 0
+ em = 4.1E7 ef = 0.89 lintnoi = 0
+ tnoia = 7.5E6 tnoib = 7.2E6 rnoia = 0.794
+ rnoib = 0.38 xpart = 0 cgso = {1.5674E-10/sw_func_tox_hv_ratio}
+ cgdo = {3.0674E-10/sw_func_tox_hv_ratio} cgbo = {0/sw_func_tox_hv_ratio} ckappas = 0.6
+ cf = 0 clc = 1E-7 cle = 0.6
+ dlc = -3.5995E-8 dwc = 0 vfbcv = -1
+ noff = 4 voffcv = -0.2104 acde = 0.4176
+ moin = 15 cgsl = {4.49025E-11/sw_func_tox_hv_ratio} cgdl = {4.49025E-11/sw_func_tox_hv_ratio}
+ ijthsrev = 0.1 ijthsfwd = 0.1 xjbvs = 1
+ bvs = 12.636 jss = 3.75E-4 jsws = 5.84E-11
+ cjs = {8.310E-04*sw_func_nsd_pw_cj} mjs = 0.295 mjsws = 0.037586
+ cjsws = {8.643094E-11*sw_func_nsd_pw_cj} cjswgs = {5.47776E-11*sw_func_nsd_pw_cj} mjswgs = 0.78692
+ pbs = 0.72468 pbsws = 0.29067 pbswgs = 0.54958
+ tnom = 30 ute = -1.4324 kt1 = -0.37073
+ kt1l = 0 kt2 = -0.019151 ua1 = 2.0117E-9
+ ub1 = -2.9862E-18 uc1 = -5.9821E-11 at = 2.9E4
+ prt = 0 njs = 1.0773 xtis = 0.76
+ tpb = 1.344E-3 tpbsw = 9.9005E-4 tpbswg = 0
+ tcj = 6.7434E-4 tcjsw = 2.493E-4 tcjswg = 0
+ tvoff = 0 saref = 2.8E-7 sbref = 1.585E-6
+ wlod = 0 ku0 = -9.9E-8 kvsat = 0.3
+ kvth0 = 1.7057E-8 tku0 = 0 llodku0 = 1
+ wlodku0 = 1 llodvth = 1 wlodvth = 1
+ lku0 = 9.6975E-7 wku0 = 2E-7 pku0 = 0
+ lkvth0 = 2.2691E-7 wkvth0 = 2.3093E-6 pkvth0 = 0
+ stk2 = 0 lodk2 = 1 steta0 = 0
+ lodeta0 = 1

.model nvhv_model_base.4 nmos
+ level = 54 lmin = 7E-7 lmax = 2.2E-6 wmin = 5E-5
+ wmax = 6E-5 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 1 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 1.16E-8
+ toxm = 1.16E-8 xj = 1.5E-7 ndep = 1.7E17
+ ngate = 1E23 nsd = 1E20 rsh = {sw_rnw}
+ rshg = 0.1 phin = 0 wint = {2.1346E-8+sw_activecd}
+ wl = 0 wln = 1 ww = 0
+ wwn = 1 wwl = 0 lint = {7.6507E-8-sw_polycd}
+ ll = 0 lln = 1 lw = 0
+ lwn = 1 lwl = 0 llc = 0
+ lwc = 0 lwlc = 0 wlc = 0
+ wwc = 0 wwlc = 0 dwg = -4.1292E-9
+ dwb = -1.6944E-9 xl = 0 xw = 0
+ dmcg = 0 dmdg = 0 dmcgt = 0
+ xgw = 0 xgl = 0 ngcon = 1
+ vth0 = 0.800438 lvth0 = -1.075632E-8 k1 = 0.923559
+ lk1 = -5.358753E-8 k2 = -4.92657E-2 lk2 = 1.037563E-8
+ k3 = -0.884 k3b = 0.43 w0 = 0
+ lpe0 = 0 lpeb = -2.182E-7 vbm = -3
+ dvtp0 = 0 dvtp1 = 0 dvt0 = 0
+ dvt1 = 0.53 dvt2 = -0.19251 dvt0w = 0.16
+ dvt1w = 6.9091E6 dvt2w = -0.036016 u0 = 3.39297E-2
+ lu0 = 3.059095E-9 ua = -9.595287E-10 lua = 2.127901E-15
+ ub = 2.645044E-18 lub = -1.032794E-24 uc = 7.074156E-11
+ luc = -2.045873E-17 ud = 0 up = 0
+ lp = 1 eu = 1.67 vsat = 1.104359E5
+ lvsat = -2.02362E-2 a0 = 0.141473 la0 = 3.245035E-7
+ ags = -0.198265 lags = 6.786261E-7 b0 = 3.2933E-8
+ b1 = 0 keta = 1.43127E-3 lketa = -1.052791E-7
+ a1 = 0 a2 = 0.659726 rdsw = 724.62
+ rdswmin = 0 rdw = 1 rdwmin = 0
+ rsw = 0 rswmin = 0 prwb = 0
+ prwg = 0 wr = 1 voff = -0.20613
+ voffl = -4.257949E-7 minv = 0 nfactor = 0.83837
+ eta0 = 0.016128 etab = -0.02983 dsub = 0.504
+ cit = -8E-4 cdsc = 0 cdscb = 0
+ cdscd = 0 pclm = -7.58976E-2 lpclm = 4.940966E-7
+ pdiblc1 = 0.21098 pdiblc2 = 2E-4 pdiblcb = -0.26831
+ drout = 0.36652 pscbe1 = 9.3731E8 pscbe2 = 1.68E-6
+ pvag = 1.99 delta = -4.586293E-4 ldelta = 2.985794E-9
+ fprout = 10.125 pdits = 0 pditsl = 0
+ pditsd = 0 vtl = 0 xn = 3
+ alpha0 = -1.062595E-5 lalpha0 = 2.237443E-11 alpha1 = 0.573481
+ lalpha1 = 2.99923E-7 beta0 = 24.125575 lbeta0 = 2.78276E-5
+ aigbacc = 1 bigbacc = 0 cigbacc = 0
+ nigbacc = 1 aigbinv = 0.35 bigbinv = 0.03
+ cigbinv = 6E-3 eigbinv = 1.1 nigbinv = 3
+ aigc = 0.43 bigc = 0.054 cigc = 0.075
+ aigsd = 0.43 bigsd = 0.054 cigsd = 0.075
+ dlcig = 0 nigc = 1 poxedge = 1
+ pigcd = 1 ntox = 1 toxref = 1.16E-8
+ agidl = 0 bgidl = 1.058E9 cgidl = 4E3
+ egidl = 0.8 noia = 2.6E41 noib = 0
+ noic = 0 em = 4.1E7 ef = 0.89
+ lintnoi = 0 tnoia = 7.5E6 tnoib = 7.2E6
+ rnoia = 0.794 rnoib = 0.38 xpart = 0
+ cgso = {1.5674E-10/sw_func_tox_hv_ratio} cgdo = {3.0674E-10/sw_func_tox_hv_ratio} cgbo = {0/sw_func_tox_hv_ratio}
+ ckappas = 0.6 cf = 0 clc = 1E-7
+ cle = 0.6 dlc = -3.5995E-8 dwc = 0
+ vfbcv = -1 noff = 4 voffcv = -0.2104
+ acde = 0.4176 moin = 15 cgsl = {4.49025E-11/sw_func_tox_hv_ratio}
+ cgdl = {4.49025E-11/sw_func_tox_hv_ratio} ijthsrev = 0.1 ijthsfwd = 0.1
+ xjbvs = 1 bvs = 12.636 jss = 3.75E-4
+ jsws = 5.84E-11 cjs = {8.310E-04*sw_func_nsd_pw_cj} mjs = 0.295
+ mjsws = 0.037586 cjsws = {8.643094E-11*sw_func_nsd_pw_cj} cjswgs = {5.47776E-11*sw_func_nsd_pw_cj}
+ mjswgs = 0.78692 pbs = 0.72468 pbsws = 0.29067
+ pbswgs = 0.54958 tnom = 30 ute = -1.417741
+ lute = -3.000723E-8 kt1 = -0.37073 kt1l = 0
+ kt2 = -3.181197E-3 lkt2 = -3.268996E-8 ua1 = 2.0117E-9
+ ub1 = -3.237121E-18 lub1 = 5.136312E-25 uc1 = -8.080006E-11
+ luc1 = 4.294385E-17 at = 2.9E4 prt = 0
+ njs = 1.0773 xtis = 0.76 tpb = 1.344E-3
+ tpbsw = 9.9005E-4 tpbswg = 0 tcj = 6.7434E-4
+ tcjsw = 2.493E-4 tcjswg = 0 tvoff = 0
+ saref = 2.8E-7 sbref = 1.585E-6 wlod = 0
+ ku0 = -9.9E-8 kvsat = 0.3 kvth0 = 1.7057E-8
+ tku0 = 0 llodku0 = 1 wlodku0 = 1
+ llodvth = 1 wlodvth = 1 lku0 = 9.6975E-7
+ wku0 = 2E-7 pku0 = 0 lkvth0 = 2.2691E-7
+ wkvth0 = 2.3093E-6 pkvth0 = 0 stk2 = 0
+ lodk2 = 1 steta0 = 0 lodeta0 = 1

.model nvhv_model_base.5 nmos
+ level = 54 lmin = 2.2E-6 lmax = 2.02E-5 wmin = 2E-5
+ wmax = 5E-5 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 1 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 1.16E-8
+ toxm = 1.16E-8 xj = 1.5E-7 ndep = 1.7E17
+ ngate = 1E23 nsd = 1E20 rsh = {sw_rnw}
+ rshg = 0.1 phin = 0 wint = {2.1346E-8+sw_activecd}
+ wl = 0 wln = 1 ww = 0
+ wwn = 1 wwl = 0 lint = {7.6507E-8-sw_polycd}
+ ll = 0 lln = 1 lw = 0
+ lwn = 1 lwl = 0 llc = 0
+ lwc = 0 lwlc = 0 wlc = 0
+ wwc = 0 wwlc = 0 dwg = -4.1292E-9
+ dwb = -1.6944E-9 xl = 0 xw = 0
+ dmcg = 0 dmdg = 0 dmcgt = 0
+ xgw = 0 xgl = 0 ngcon = 1
+ vth0 = 0.795183 k1 = 0.89738 k2 = -0.044197
+ k3 = -0.884 k3b = 0.43 w0 = 0
+ lpe0 = 0 lpeb = -2.182E-7 vbm = -3
+ dvtp0 = 0 dvtp1 = 0 dvt0 = 0
+ dvt1 = 0.53 dvt2 = -0.19251 dvt0w = 0.16
+ dvt1w = 6.9091E6 dvt2w = -0.036016 u0 = 3.54241E-2
+ ua = 8E-11 ub = 2.1405E-18 uc = 6.0747E-11
+ ud = 0 up = 0 lp = 1
+ eu = 1.67 vsat = 1.0055E5 a0 = 0.3
+ ags = 0.13326 b0 = 3.2933E-8 b1 = 0
+ keta = -0.05 a1 = 0 a2 = 0.659726
+ rdsw = 724.62 rdswmin = 0 rdw = 1
+ rdwmin = 0 rsw = 0 rswmin = 0
+ prwb = 0 prwg = 0 wr = 1
+ voff = -0.20613 voffl = -4.257949E-7 minv = 0
+ nfactor = 0.83837 eta0 = 0.016128 etab = -0.02983
+ dsub = 0.504 cit = -8E-4 cdsc = 0
+ cdscb = 0 cdscd = 0 pclm = 0.16548
+ pdiblc1 = 0.21098 pdiblc2 = 2E-4 pdiblcb = -0.26831
+ drout = 0.36652 pscbe1 = 9.3731E8 pscbe2 = 1.68E-6
+ pvag = 1.99 delta = 1E-3 fprout = 10.125
+ pdits = 0 pditsl = 0 pditsd = 0
+ vtl = 0 xn = 3 alpha0 = 3.0448E-7
+ alpha1 = 0.72 beta0 = 37.72 aigbacc = 1
+ bigbacc = 0 cigbacc = 0 nigbacc = 1
+ aigbinv = 0.35 bigbinv = 0.03 cigbinv = 6E-3
+ eigbinv = 1.1 nigbinv = 3 aigc = 0.43
+ bigc = 0.054 cigc = 0.075 aigsd = 0.43
+ bigsd = 0.054 cigsd = 0.075 dlcig = 0
+ nigc = 1 poxedge = 1 pigcd = 1
+ ntox = 1 toxref = 1.16E-8 agidl = 0
+ bgidl = 1.058E9 cgidl = 4E3 egidl = 0.8
+ noia = 2.6E41 noib = 0 noic = 0
+ em = 4.1E7 ef = 0.89 lintnoi = 0
+ tnoia = 7.5E6 tnoib = 7.2E6 rnoia = 0.794
+ rnoib = 0.38 xpart = 0 cgso = {1.5674E-10/sw_func_tox_hv_ratio}
+ cgdo = {3.0674E-10/sw_func_tox_hv_ratio} cgbo = {0/sw_func_tox_hv_ratio} ckappas = 0.6
+ cf = 0 clc = 1E-7 cle = 0.6
+ dlc = -3.5995E-8 dwc = 0 vfbcv = -1
+ noff = 4 voffcv = -0.2104 acde = 0.4176
+ moin = 15 cgsl = {4.49025E-11/sw_func_tox_hv_ratio} cgdl = {4.49025E-11/sw_func_tox_hv_ratio}
+ ijthsrev = 0.1 ijthsfwd = 0.1 xjbvs = 1
+ bvs = 12.636 jss = 3.75E-4 jsws = 5.84E-11
+ cjs = {8.310E-04*sw_func_nsd_pw_cj} mjs = 0.295 mjsws = 0.037586
+ cjsws = {8.643094E-11*sw_func_nsd_pw_cj} cjswgs = {5.47776E-11*sw_func_nsd_pw_cj} mjswgs = 0.78692
+ pbs = 0.72468 pbsws = 0.29067 pbswgs = 0.54958
+ tnom = 30 ute = -1.4324 kt1 = -0.37073
+ kt1l = 0 kt2 = -0.019151 ua1 = 2.0117E-9
+ ub1 = -2.9862E-18 uc1 = -5.9821E-11 at = 2.9E4
+ prt = 0 njs = 1.0773 xtis = 0.76
+ tpb = 1.344E-3 tpbsw = 9.9005E-4 tpbswg = 0
+ tcj = 6.7434E-4 tcjsw = 2.493E-4 tcjswg = 0
+ tvoff = 0 saref = 2.8E-7 sbref = 1.585E-6
+ wlod = 0 ku0 = -9.9E-8 kvsat = 0.3
+ kvth0 = 1.7057E-8 tku0 = 0 llodku0 = 1
+ wlodku0 = 1 llodvth = 1 wlodvth = 1
+ lku0 = 9.6975E-7 wku0 = 2E-7 pku0 = 0
+ lkvth0 = 2.2691E-7 wkvth0 = 2.3093E-6 pkvth0 = 0
+ stk2 = 0 lodk2 = 1 steta0 = 0
+ lodeta0 = 1

.model nvhv_model_base.6 nmos
+ level = 54 lmin = 7E-7 lmax = 2.2E-6 wmin = 2E-5
+ wmax = 5E-5 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 1 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 1.16E-8
+ toxm = 1.16E-8 xj = 1.5E-7 ndep = 1.7E17
+ ngate = 1E23 nsd = 1E20 rsh = {sw_rnw}
+ rshg = 0.1 phin = 0 wint = {2.1346E-8+sw_activecd}
+ wl = 0 wln = 1 ww = 0
+ wwn = 1 wwl = 0 lint = {7.6507E-8-sw_polycd}
+ ll = 0 lln = 1 lw = 0
+ lwn = 1 lwl = 0 llc = 0
+ lwc = 0 lwlc = 0 wlc = 0
+ wwc = 0 wwlc = 0 dwg = -4.1292E-9
+ dwb = -1.6944E-9 xl = 0 xw = 0
+ dmcg = 0 dmdg = 0 dmcgt = 0
+ xgw = 0 xgl = 0 ngcon = 1
+ vth0 = 0.800901 lvth0 = -1.170378E-8 wvth0 = -2.312294E-8
+ pvth0 = 4.733233E-14 k1 = 0.923559 lk1 = -5.358753E-8
+ k2 = -4.91942E-2 lk2 = 1.022915E-8 wk2 = -3.575088E-9
+ pk2 = 7.318154E-15 k3 = -0.884 k3b = 0.43
+ w0 = 0 lpe0 = 0 lpeb = -2.182E-7
+ vbm = -3 dvtp0 = 0 dvtp1 = 0
+ dvt0 = 0 dvt1 = 0.53 dvt2 = -0.19251
+ dvt0w = 0.16 dvt1w = 6.9091E6 dvt2w = -0.036016
+ u0 = 3.40302E-2 lu0 = 2.853366E-9 wu0 = -5.020877E-9
+ pu0 = 1.027767E-14 ua = -1.097123E-9 lua = 2.409555E-15
+ wua = 6.873864E-15 pua = -1.40707E-20 ub = 2.737423E-18
+ lub = -1.221892E-24 wub = -4.615014E-24 pub = 9.446869E-30
+ uc = 6.809037E-11 luc = -1.503177E-17 wuc = 1.324467E-16
+ puc = -2.711165E-22 ud = 0 up = 0
+ lp = 1 eu = 1.67 vsat = 1.104359E5
+ lvsat = -2.02362E-2 a0 = 0.141473 la0 = 3.245035E-7
+ ags = -0.198265 lags = 6.786261E-7 b0 = 3.2933E-8
+ b1 = 0 keta = 1.43127E-3 lketa = -1.052791E-7
+ a1 = 0 a2 = 0.659726 rdsw = 724.62
+ rdswmin = 0 rdw = 1 rdwmin = 0
+ rsw = 0 rswmin = 0 prwb = 0
+ prwg = 0 wr = 1 voff = -0.20613
+ voffl = -4.257949E-7 minv = 0 nfactor = 0.83837
+ eta0 = 0.016128 etab = -0.02983 dsub = 0.504
+ cit = -8E-4 cdsc = 0 cdscb = 0
+ cdscd = 0 pclm = -7.58976E-2 lpclm = 4.940966E-7
+ pdiblc1 = 0.21098 pdiblc2 = 2E-4 pdiblcb = -0.26831
+ drout = 0.36652 pscbe1 = 9.3731E8 pscbe2 = 1.68E-6
+ pvag = 1.99 delta = -4.586293E-4 ldelta = 2.985794E-9
+ fprout = 10.125 pdits = 0 pditsl = 0
+ pditsd = 0 vtl = 0 xn = 3
+ alpha0 = -1.062595E-5 lalpha0 = 2.237443E-11 alpha1 = 0.573481
+ lalpha1 = 2.99923E-7 beta0 = 24.125575 lbeta0 = 2.78276E-5
+ aigbacc = 1 bigbacc = 0 cigbacc = 0
+ nigbacc = 1 aigbinv = 0.35 bigbinv = 0.03
+ cigbinv = 6E-3 eigbinv = 1.1 nigbinv = 3
+ aigc = 0.43 bigc = 0.054 cigc = 0.075
+ aigsd = 0.43 bigsd = 0.054 cigsd = 0.075
+ dlcig = 0 nigc = 1 poxedge = 1
+ pigcd = 1 ntox = 1 toxref = 1.16E-8
+ agidl = 0 bgidl = 1.058E9 cgidl = 4E3
+ egidl = 0.8 noia = 2.6E41 noib = 0
+ noic = 0 em = 4.1E7 ef = 0.89
+ lintnoi = 0 tnoia = 7.5E6 tnoib = 7.2E6
+ rnoia = 0.794 rnoib = 0.38 xpart = 0
+ cgso = {1.5674E-10/sw_func_tox_hv_ratio} cgdo = {3.0674E-10/sw_func_tox_hv_ratio} cgbo = {0/sw_func_tox_hv_ratio}
+ ckappas = 0.6 cf = 0 clc = 1E-7
+ cle = 0.6 dlc = -3.5995E-8 dwc = 0
+ vfbcv = -1 noff = 4 voffcv = -0.2104
+ acde = 0.4176 moin = 15 cgsl = {4.49025E-11/sw_func_tox_hv_ratio}
+ cgdl = {4.49025E-11/sw_func_tox_hv_ratio} ijthsrev = 0.1 ijthsfwd = 0.1
+ xjbvs = 1 bvs = 12.636 jss = 3.75E-4
+ jsws = 5.84E-11 cjs = {8.310E-04*sw_func_nsd_pw_cj} mjs = 0.295
+ mjsws = 0.037586 cjsws = {8.643094E-11*sw_func_nsd_pw_cj} cjswgs = {5.47776E-11*sw_func_nsd_pw_cj}
+ mjswgs = 0.78692 pbs = 0.72468 pbsws = 0.29067
+ pbswgs = 0.54958 tnom = 30 ute = -1.363038
+ lute = -1.419838E-7 wute = -2.732821E-6 pute = 5.594047E-12
+ kt1 = -0.37073 kt1l = 0 kt2 = 7.442613E-3
+ lkt2 = -5.443675E-8 wkt2 = -5.307369E-7 pkt2 = 1.086411E-12
+ ua1 = 2.0117E-9 ub1 = -3.237121E-18 lub1 = 5.136312E-25
+ uc1 = -9.382739E-11 luc1 = 6.961061E-17 wuc1 = 6.508102E-16
+ puc1 = -1.332199E-21 at = 2.9E4 prt = 0
+ njs = 1.0773 xtis = 0.76 tpb = 1.344E-3
+ tpbsw = 9.9005E-4 tpbswg = 0 tcj = 6.7434E-4
+ tcjsw = 2.493E-4 tcjswg = 0 tvoff = 0
+ saref = 2.8E-7 sbref = 1.585E-6 wlod = 0
+ ku0 = -9.9E-8 kvsat = 0.3 kvth0 = 1.7057E-8
+ tku0 = 0 llodku0 = 1 wlodku0 = 1
+ llodvth = 1 wlodvth = 1 lku0 = 9.6975E-7
+ wku0 = 2E-7 pku0 = 0 lkvth0 = 2.2691E-7
+ wkvth0 = 2.3093E-6 pkvth0 = 0 stk2 = 0
+ lodk2 = 1 steta0 = 0 lodeta0 = 1

.model nvhv_model_base.7 nmos
+ level = 54 lmin = 2.2E-6 lmax = 2.02E-5 wmin = 5E-6
+ wmax = 2E-5 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 1 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 1.16E-8
+ toxm = 1.16E-8 xj = 1.5E-7 ndep = 1.7E17
+ ngate = 1E23 nsd = 1E20 rsh = {sw_rnw}
+ rshg = 0.1 phin = 0 wint = {2.1346E-8+sw_activecd}
+ wl = 0 wln = 1 ww = 0
+ wwn = 1 wwl = 0 lint = {7.6507E-8-sw_polycd}
+ ll = 0 lln = 1 lw = 0
+ lwn = 1 lwl = 0 llc = 0
+ lwc = 0 lwlc = 0 wlc = 0
+ wwc = 0 wwlc = 0 dwg = -4.1292E-9
+ dwb = -1.6944E-9 xl = 0 xw = 0
+ dmcg = 0 dmdg = 0 dmcgt = 0
+ xgw = 0 xgl = 0 ngcon = 1
+ vth0 = 0.792999 wvth0 = 4.358396E-8 k1 = 0.89738
+ k2 = -0.044197 k3 = -0.884 k3b = 0.43
+ w0 = 0 lpe0 = 0 lpeb = -2.182E-7
+ vbm = -3 dvtp0 = 0 dvtp1 = 0
+ dvt0 = 0 dvt1 = 0.53 dvt2 = -0.19251
+ dvt0w = 0.16 dvt1w = 6.9091E6 dvt2w = -0.036016
+ u0 = 3.59523E-2 wu0 = -1.054114E-8 ua = 8E-11
+ ub = 2.264995E-18 wub = -2.484576E-24 uc = 7.198951E-11
+ wuc = -2.243703E-16 ud = 0 up = 0
+ lp = 1 eu = 1.67 vsat = 1.0055E5
+ a0 = 0.3 ags = 0.13326 b0 = 3.2933E-8
+ b1 = 0 keta = -0.05 a1 = 0
+ a2 = 0.659726 rdsw = 724.62 rdswmin = 0
+ rdw = 1 rdwmin = 0 rsw = 0
+ rswmin = 0 prwb = 0 prwg = 0
+ wr = 1 voff = -0.20613 voffl = -4.257949E-7
+ minv = 0 nfactor = 0.83837 eta0 = 0.016128
+ etab = -0.02983 dsub = 0.504 cit = -8E-4
+ cdsc = 0 cdscb = 0 cdscd = 0
+ pclm = 0.16548 pdiblc1 = 0.21098 pdiblc2 = 2E-4
+ pdiblcb = -0.26831 drout = 0.36652 pscbe1 = 9.3731E8
+ pscbe2 = 1.68E-6 pvag = 1.99 delta = 1E-3
+ fprout = 10.125 pdits = 0 pditsl = 0
+ pditsd = 0 vtl = 0 xn = 3
+ alpha0 = 3.0448E-7 alpha1 = 0.72 beta0 = 37.72
+ aigbacc = 1 bigbacc = 0 cigbacc = 0
+ nigbacc = 1 aigbinv = 0.35 bigbinv = 0.03
+ cigbinv = 6E-3 eigbinv = 1.1 nigbinv = 3
+ aigc = 0.43 bigc = 0.054 cigc = 0.075
+ aigsd = 0.43 bigsd = 0.054 cigsd = 0.075
+ dlcig = 0 nigc = 1 poxedge = 1
+ pigcd = 1 ntox = 1 toxref = 1.16E-8
+ agidl = 0 bgidl = 1.058E9 cgidl = 4E3
+ egidl = 0.8 noia = 2.6E41 noib = 0
+ noic = 0 em = 4.1E7 ef = 0.89
+ lintnoi = 0 tnoia = 7.5E6 tnoib = 7.2E6
+ rnoia = 0.794 rnoib = 0.38 xpart = 0
+ cgso = {1.5674E-10/sw_func_tox_hv_ratio} cgdo = {3.0674E-10/sw_func_tox_hv_ratio} cgbo = {0/sw_func_tox_hv_ratio}
+ ckappas = 0.6 cf = 0 clc = 1E-7
+ cle = 0.6 dlc = -3.5995E-8 dwc = 0
+ vfbcv = -1 noff = 4 voffcv = -0.2104
+ acde = 0.4176 moin = 15 cgsl = {4.49025E-11/sw_func_tox_hv_ratio}
+ cgdl = {4.49025E-11/sw_func_tox_hv_ratio} ijthsrev = 0.1 ijthsfwd = 0.1
+ xjbvs = 1 bvs = 12.636 jss = 3.75E-4
+ jsws = 5.84E-11 cjs = {8.310E-04*sw_func_nsd_pw_cj} mjs = 0.295
+ mjsws = 0.037586 cjsws = {8.643094E-11*sw_func_nsd_pw_cj} cjswgs = {5.47776E-11*sw_func_nsd_pw_cj}
+ mjswgs = 0.78692 pbs = 0.72468 pbsws = 0.29067
+ pbswgs = 0.54958 tnom = 30 ute = -1.4324
+ kt1 = -0.37073 kt1l = 0 kt2 = -0.019151
+ ua1 = 2.0117E-9 ub1 = -3.004476E-18 wub1 = 3.647386E-25
+ uc1 = -5.9821E-11 at = 2.9E4 prt = 0
+ njs = 1.0773 xtis = 0.76 tpb = 1.344E-3
+ tpbsw = 9.9005E-4 tpbswg = 0 tcj = 6.7434E-4
+ tcjsw = 2.493E-4 tcjswg = 0 tvoff = 0
+ saref = 2.8E-7 sbref = 1.585E-6 wlod = 0
+ ku0 = -9.9E-8 kvsat = 0.3 kvth0 = 1.7057E-8
+ tku0 = 0 llodku0 = 1 wlodku0 = 1
+ llodvth = 1 wlodvth = 1 lku0 = 9.6975E-7
+ wku0 = 2E-7 pku0 = 0 lkvth0 = 2.2691E-7
+ wkvth0 = 2.3093E-6 pkvth0 = 0 stk2 = 0
+ lodk2 = 1 steta0 = 0 lodeta0 = 1

.model nvhv_model_base.8 nmos
+ level = 54 lmin = 7E-7 lmax = 2.2E-6 wmin = 5E-6
+ wmax = 2E-5 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 1 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 1.16E-8
+ toxm = 1.16E-8 xj = 1.5E-7 ndep = 1.7E17
+ ngate = 1E23 nsd = 1E20 rsh = {sw_rnw}
+ rshg = 0.1 phin = 0 wint = {2.1346E-8+sw_activecd}
+ wl = 0 wln = 1 ww = 0
+ wwn = 1 wwl = 0 lint = {7.6507E-8-sw_polycd}
+ ll = 0 lln = 1 lw = 0
+ lwn = 1 lwl = 0 llc = 0
+ lwc = 0 lwlc = 0 wlc = 0
+ wwc = 0 wwlc = 0 dwg = -4.1292E-9
+ dwb = -1.6944E-9 xl = 0 xw = 0
+ dmcg = 0 dmdg = 0 dmcgt = 0
+ xgw = 0 xgl = 0 ngcon = 1
+ vth0 = 0.797079 lvth0 = -8.351253E-9 wvth0 = 5.314682E-8
+ pvth0 = -1.957505E-14 k1 = 0.93221 lk1 = -7.129753E-8
+ wk1 = -1.726655E-7 pk1 = 3.534438E-13 k2 = -5.14456E-2
+ lk2 = 1.48377E-8 wk2 = 4.13565E-8 pk2 = -8.465617E-14
+ k3 = -0.884 k3b = 0.43 w0 = 0
+ lpe0 = 0 lpeb = -2.182E-7 vbm = -3
+ dvtp0 = 0 dvtp1 = 0 dvt0 = 0
+ dvt1 = 0.53 dvt2 = -0.19251 dvt0w = 0.16
+ dvt1w = 6.9091E6 dvt2w = -0.036016 u0 = 3.32905E-2
+ lu0 = 5.448576E-9 wu0 = 9.740255E-9 pu0 = -4.151574E-14
+ ua = -9.550993E-10 lua = 2.118834E-15 wua = 4.039444E-15
+ pua = -8.268685E-21 ub = 2.72512E-18 lub = -9.418708E-25
+ wub = -4.369489E-24 pub = 3.858391E-30 uc = 8.547057E-11
+ luc = -2.759554E-17 wuc = -2.144154E-16 puc = -2.037754E-23
+ ud = 0 up = 0 lp = 1
+ eu = 1.67 vsat = 1.104359E5 lvsat = -2.02362E-2
+ a0 = 0.141473 la0 = 3.245035E-7 ags = -0.198265
+ lags = 6.786261E-7 b0 = 3.2933E-8 b1 = 0
+ keta = 1.43127E-3 lketa = -1.052791E-7 a1 = 0
+ a2 = 0.659726 rdsw = 724.62 rdswmin = 0
+ rdw = 1 rdwmin = 0 rsw = 0
+ rswmin = 0 prwb = 0 prwg = 0
+ wr = 1 voff = -0.20613 voffl = -4.257949E-7
+ minv = 0 nfactor = 0.83837 eta0 = 0.016128
+ etab = -0.02983 dsub = 0.504 cit = -8E-4
+ cdsc = 0 cdscb = 0 cdscd = 0
+ pclm = -7.58976E-2 lpclm = 4.940966E-7 pdiblc1 = 0.21098
+ pdiblc2 = 2E-4 pdiblcb = -0.26831 drout = 0.36652
+ pscbe1 = 9.3731E8 pscbe2 = 1.68E-6 pvag = 1.99
+ delta = -4.586293E-4 ldelta = 2.985794E-9 fprout = 10.125
+ pdits = 0 pditsl = 0 pditsd = 0
+ vtl = 0 xn = 3 alpha0 = -1.062595E-5
+ lalpha0 = 2.237443E-11 alpha1 = 0.573481 lalpha1 = 2.99923E-7
+ beta0 = 24.125575 lbeta0 = 2.78276E-5 aigbacc = 1
+ bigbacc = 0 cigbacc = 0 nigbacc = 1
+ aigbinv = 0.35 bigbinv = 0.03 cigbinv = 6E-3
+ eigbinv = 1.1 nigbinv = 3 aigc = 0.43
+ bigc = 0.054 cigc = 0.075 aigsd = 0.43
+ bigsd = 0.054 cigsd = 0.075 dlcig = 0
+ nigc = 1 poxedge = 1 pigcd = 1
+ ntox = 1 toxref = 1.16E-8 agidl = 0
+ bgidl = 1.058E9 cgidl = 4E3 egidl = 0.8
+ noia = 2.6E41 noib = 0 noic = 0
+ em = 4.1E7 ef = 0.89 lintnoi = 0
+ tnoia = 7.5E6 tnoib = 7.2E6 rnoia = 0.794
+ rnoib = 0.38 xpart = 0 cgso = {1.5674E-10/sw_func_tox_hv_ratio}
+ cgdo = {3.0674E-10/sw_func_tox_hv_ratio} cgbo = {0/sw_func_tox_hv_ratio} ckappas = 0.6
+ cf = 0 clc = 1E-7 cle = 0.6
+ dlc = -3.5995E-8 dwc = 0 vfbcv = -1
+ noff = 4 voffcv = -0.2104 acde = 0.4176
+ moin = 15 cgsl = {4.49025E-11/sw_func_tox_hv_ratio} cgdl = {4.49025E-11/sw_func_tox_hv_ratio}
+ ijthsrev = 0.1 ijthsfwd = 0.1 xjbvs = 1
+ bvs = 12.636 jss = 3.75E-4 jsws = 5.84E-11
+ cjs = {8.310E-04*sw_func_nsd_pw_cj} mjs = 0.295 mjsws = 0.037586
+ cjsws = {8.643094E-11*sw_func_nsd_pw_cj} cjswgs = {5.47776E-11*sw_func_nsd_pw_cj} mjswgs = 0.78692
+ pbs = 0.72468 pbsws = 0.29067 pbswgs = 0.54958
+ tnom = 30 ute = -1.499971 lute = 1.383169E-7
+ kt1 = -0.37073 kt1l = 0 kt2 = -0.019151
+ ua1 = 2.0117E-9 ub1 = -3.262061E-18 lub1 = 5.272732E-25
+ wub1 = 4.977432E-25 pub1 = -2.722586E-31 uc1 = -6.167872E-11
+ luc1 = 3.802734E-18 wuc1 = 9.209306E-18 puc1 = -1.885132E-23
+ at = 2.9E4 prt = 0 njs = 1.0773
+ xtis = 0.76 tpb = 1.344E-3 tpbsw = 9.9005E-4
+ tpbswg = 0 tcj = 6.7434E-4 tcjsw = 2.493E-4
+ tcjswg = 0 tvoff = 0 saref = 2.8E-7
+ sbref = 1.585E-6 wlod = 0 ku0 = -9.9E-8
+ kvsat = 0.3 kvth0 = 1.7057E-8 tku0 = 0
+ llodku0 = 1 wlodku0 = 1 llodvth = 1
+ wlodvth = 1 lku0 = 9.6975E-7 wku0 = 2E-7
+ pku0 = 0 lkvth0 = 2.2691E-7 wkvth0 = 2.3093E-6
+ pkvth0 = 0 stk2 = 0 lodk2 = 1
+ steta0 = 0 lodeta0 = 1

.ends sky130_fd_pr__nfet_g5v0d16v0_base
