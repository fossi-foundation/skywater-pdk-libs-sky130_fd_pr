library sky130.lib

// * Copyright 2022 The SkyWater PDK Authors
section tt
parameters mc_mm_switch=0
parameters mc_pr_switch=0
parameters corner_factor=1
parameters process_mc_factor=1
parameters mismatch_factor=1
include "continuous/parameters_fet_tt.scs"
include "continuous/parameters_res_nom.scs"
include "continuous/parameters_cap_nom.scs"
include "continuous/models_global.scs"
include "continuous/models_fet.scs"
include "continuous/models_bjt.scs"
include "continuous/models_diodes.scs"
include "continuous/models_resistors.scs"
include "continuous/models_capacitors.scs"
include "corners/tt.scs"
include "corners/tt/specialized_cells.scs"
include "rescap/res_typical__cap_typical.scs"
include "rescap/res_typical__cap_typical__lin.scs"
endsection tt

section sf
parameters mc_mm_switch=0
parameters mc_pr_switch=0
parameters corner_factor=1
parameters process_mc_factor=1
parameters mismatch_factor=1
include "continuous/parameters_fet_sf.scs"
include "continuous/parameters_res_nom.scs"
include "continuous/parameters_cap_nom.scs"
include "continuous/models_global.scs"
include "continuous/models_fet.scs"
include "continuous/models_bjt.scs"
include "continuous/models_diodes.scs"
include "continuous/models_resistors.scs"
include "continuous/models_capacitors.scs"
include "corners/sf.scs"
include "corners/sf/specialized_cells.scs"
include "rescap/res_typical__cap_typical.scs"
include "rescap/res_typical__cap_typical__lin.scs"
endsection sf

section ff
parameters mc_mm_switch=0
parameters mc_pr_switch=0
parameters corner_factor=1
parameters process_mc_factor=1
parameters mismatch_factor=1
include "continuous/parameters_fet_ff.scs"
include "continuous/parameters_res_nom.scs"
include "continuous/parameters_cap_nom.scs"
include "continuous/models_global.scs"
include "continuous/models_fet.scs"
include "continuous/models_bjt.scs"
include "continuous/models_diodes.scs"
include "continuous/models_resistors.scs"
include "continuous/models_capacitors.scs"
include "corners/ff.scs"
include "corners/ff/specialized_cells.scs"
include "rescap/res_typical__cap_typical.scs"
include "rescap/res_typical__cap_typical__lin.scs"
endsection ff

section ss
parameters mc_mm_switch=0
parameters mc_pr_switch=0
parameters corner_factor=1
parameters process_mc_factor=1
parameters mismatch_factor=1
include "continuous/parameters_fet_ss.scs"
include "continuous/parameters_res_nom.scs"
include "continuous/parameters_cap_nom.scs"
include "continuous/models_global.scs"
include "continuous/models_fet.scs"
include "continuous/models_bjt.scs"
include "continuous/models_diodes.scs"
include "continuous/models_resistors.scs"
include "continuous/models_capacitors.scs"
include "corners/ss.scs"
include "corners/ss/specialized_cells.scs"
include "rescap/res_typical__cap_typical.scs"
include "rescap/res_typical__cap_typical__lin.scs"
endsection ss

section fs
parameters mc_mm_switch=0
parameters mc_pr_switch=0
parameters corner_factor=1
parameters process_mc_factor=1
parameters mismatch_factor=1
include "continuous/parameters_fet_fs.scs"
include "continuous/parameters_res_nom.scs"
include "continuous/parameters_cap_nom.scs"
include "continuous/models_global.scs"
include "continuous/models_fet.scs"
include "continuous/models_bjt.scs"
include "continuous/models_diodes.scs"
include "continuous/models_resistors.scs"
include "continuous/models_capacitors.scs"
include "corners/fs.scs"
include "corners/fs/specialized_cells.scs"
include "rescap/res_typical__cap_typical.scs"
include "rescap/res_typical__cap_typical__lin.scs"
endsection fs

section ll
parameters mc_mm_switch=0
parameters mc_pr_switch=0
parameters corner_factor=1
parameters process_mc_factor=1
parameters mismatch_factor=1
include "continuous/parameters_fet_tt.scs"
include "continuous/parameters_res_low.scs"
include "continuous/parameters_cap_low.scs"
include "continuous/models_global.scs"
include "continuous/models_fet.scs"
include "continuous/models_bjt.scs"
include "continuous/models_diodes.scs"
include "continuous/models_resistors.scs"
include "continuous/models_capacitors.scs"
include "corners/tt.scs"
include "corners/tt/specialized_cells.scs"
include "rescap/res_low__cap_low.scs"
include "rescap/res_low__cap_low__lin.scs"
endsection ll

section hh
parameters mc_mm_switch=0
parameters mc_pr_switch=0
parameters corner_factor=1
parameters process_mc_factor=1
parameters mismatch_factor=1
include "continuous/parameters_fet_tt.scs"
include "continuous/parameters_res_high.scs"
include "continuous/parameters_cap_high.scs"
include "continuous/models_global.scs"
include "continuous/models_fet.scs"
include "continuous/models_bjt.scs"
include "continuous/models_diodes.scs"
include "continuous/models_resistors.scs"
include "continuous/models_capacitors.scs"
include "corners/tt.scs"
include "corners/tt/specialized_cells.scs"
include "rescap/res_high__cap_high.scs"
include "rescap/res_high__cap_high__lin.scs"
endsection hh

section hl
parameters mc_mm_switch=0
parameters mc_pr_switch=0
parameters corner_factor=1
parameters process_mc_factor=1
parameters mismatch_factor=1
include "continuous/parameters_fet_tt.scs"
include "continuous/parameters_res_high.scs"
include "continuous/parameters_cap_low.scs"
include "continuous/models_global.scs"
include "continuous/models_fet.scs"
include "continuous/models_bjt.scs"
include "continuous/models_diodes.scs"
include "continuous/models_resistors.scs"
include "continuous/models_capacitors.scs"
include "corners/tt.scs"
include "corners/tt/specialized_cells.scs"
include "rescap/res_high__cap_low.scs"
include "rescap/res_high__cap_low__lin.scs"
endsection hl

section lh
parameters mc_mm_switch=0
parameters mc_pr_switch=0
parameters corner_factor=1
parameters process_mc_factor=1
parameters mismatch_factor=1
include "continuous/parameters_fet_tt.scs"
include "continuous/parameters_res_low.scs"
include "continuous/parameters_cap_high.scs"
include "continuous/models_global.scs"
include "continuous/models_fet.scs"
include "continuous/models_bjt.scs"
include "continuous/models_diodes.scs"
include "continuous/models_resistors.scs"
include "continuous/models_capacitors.scs"
include "corners/tt.scs"
include "corners/tt/specialized_cells.scs"
include "rescap/res_low__cap_high.scs"
include "rescap/res_low__cap_high__lin.scs"
endsection lh

section ss_ll
parameters mc_mm_switch=0
parameters mc_pr_switch=0
parameters corner_factor=1
parameters process_mc_factor=1
parameters mismatch_factor=1
include "continuous/parameters_fet_ss.scs"
include "continuous/parameters_res_low.scs"
include "continuous/parameters_cap_low.scs"
include "continuous/models_global.scs"
include "continuous/models_fet.scs"
include "continuous/models_bjt.scs"
include "continuous/models_diodes.scs"
include "continuous/models_resistors.scs"
include "continuous/models_capacitors.scs"
include "corners/ss.scs"
include "corners/ss/specialized_cells.scs"
include "rescap/res_low__cap_low.scs"
include "rescap/res_low__cap_low__lin.scs"
endsection ss_ll

section ss_hl
parameters mc_mm_switch=0
parameters mc_pr_switch=0
parameters corner_factor=1
parameters process_mc_factor=1
parameters mismatch_factor=1
include "continuous/parameters_fet_ss.scs"
include "continuous/parameters_res_high.scs"
include "continuous/parameters_cap_low.scs"
include "continuous/models_global.scs"
include "continuous/models_fet.scs"
include "continuous/models_bjt.scs"
include "continuous/models_diodes.scs"
include "continuous/models_resistors.scs"
include "continuous/models_capacitors.scs"
include "corners/ss.scs"
include "corners/ss/specialized_cells.scs"
include "rescap/res_high__cap_low.scs"
include "rescap/res_high__cap_low__lin.scs"
endsection ss_hl

section ss_lh
parameters mc_mm_switch=0
parameters mc_pr_switch=0
parameters corner_factor=1
parameters process_mc_factor=1
parameters mismatch_factor=1
include "continuous/parameters_fet_ss.scs"
include "continuous/parameters_res_low.scs"
include "continuous/parameters_cap_high.scs"
include "continuous/models_global.scs"
include "continuous/models_fet.scs"
include "continuous/models_bjt.scs"
include "continuous/models_diodes.scs"
include "continuous/models_resistors.scs"
include "continuous/models_capacitors.scs"
include "corners/ss.scs"
include "corners/ss/specialized_cells.scs"
include "rescap/res_low__cap_high.scs"
include "rescap/res_low__cap_high__lin.scs"
endsection ss_lh

section ss_hh
parameters mc_mm_switch=0
parameters mc_pr_switch=0
parameters corner_factor=1
parameters process_mc_factor=1
parameters mismatch_factor=1
include "continuous/parameters_fet_ss.scs"
include "continuous/parameters_res_high.scs"
include "continuous/parameters_cap_high.scs"
include "continuous/models_global.scs"
include "continuous/models_fet.scs"
include "continuous/models_bjt.scs"
include "continuous/models_diodes.scs"
include "continuous/models_resistors.scs"
include "continuous/models_capacitors.scs"
include "corners/ss.scs"
include "corners/ss/specialized_cells.scs"
include "rescap/res_high__cap_high.scs"
include "rescap/res_high__cap_high__lin.scs"
endsection ss_hh

section sf_ll
parameters mc_mm_switch=0
parameters mc_pr_switch=0
parameters corner_factor=1
parameters process_mc_factor=1
parameters mismatch_factor=1
include "continuous/parameters_fet_sf.scs"
include "continuous/parameters_res_low.scs"
include "continuous/parameters_cap_low.scs"
include "continuous/models_global.scs"
include "continuous/models_fet.scs"
include "continuous/models_bjt.scs"
include "continuous/models_diodes.scs"
include "continuous/models_resistors.scs"
include "continuous/models_capacitors.scs"
include "corners/sf.scs"
include "corners/sf/specialized_cells.scs"
include "rescap/res_low__cap_low.scs"
include "rescap/res_low__cap_low__lin.scs"
endsection sf_ll

section sf_hl
parameters mc_mm_switch=0
parameters mc_pr_switch=0
parameters corner_factor=1
parameters process_mc_factor=1
parameters mismatch_factor=1
include "continuous/parameters_fet_sf.scs"
include "continuous/parameters_res_high.scs"
include "continuous/parameters_cap_low.scs"
include "continuous/models_global.scs"
include "continuous/models_fet.scs"
include "continuous/models_bjt.scs"
include "continuous/models_diodes.scs"
include "continuous/models_resistors.scs"
include "continuous/models_capacitors.scs"
include "corners/sf.scs"
include "corners/sf/specialized_cells.scs"
include "rescap/res_high__cap_low.scs"
include "rescap/res_high__cap_low__lin.scs"
endsection sf_hl

section sf_hh
parameters mc_mm_switch=0
parameters mc_pr_switch=0
parameters corner_factor=1
parameters process_mc_factor=1
parameters mismatch_factor=1
include "continuous/parameters_fet_sf.scs"
include "continuous/parameters_res_high.scs"
include "continuous/parameters_cap_high.scs"
include "continuous/models_global.scs"
include "continuous/models_fet.scs"
include "continuous/models_bjt.scs"
include "continuous/models_diodes.scs"
include "continuous/models_resistors.scs"
include "continuous/models_capacitors.scs"
include "corners/sf.scs"
include "corners/sf/specialized_cells.scs"
include "rescap/res_high__cap_high.scs"
include "rescap/res_high__cap_high__lin.scs"
endsection sf_hh

section fs_ll
parameters mc_mm_switch=0
parameters mc_pr_switch=0
parameters corner_factor=1
parameters process_mc_factor=1
parameters mismatch_factor=1
include "continuous/parameters_fet_fs.scs"
include "continuous/parameters_res_low.scs"
include "continuous/parameters_cap_low.scs"
include "continuous/models_global.scs"
include "continuous/models_fet.scs"
include "continuous/models_bjt.scs"
include "continuous/models_diodes.scs"
include "continuous/models_resistors.scs"
include "continuous/models_capacitors.scs"
include "corners/fs.scs"
include "corners/fs/specialized_cells.scs"
include "rescap/res_low__cap_low.scs"
include "rescap/res_low__cap_low__lin.scs"
endsection fs_ll

section fs_hl
parameters mc_mm_switch=0
parameters mc_pr_switch=0
parameters corner_factor=1
parameters process_mc_factor=1
parameters mismatch_factor=1
include "continuous/parameters_fet_fs.scs"
include "continuous/parameters_res_high.scs"
include "continuous/parameters_cap_low.scs"
include "continuous/models_global.scs"
include "continuous/models_fet.scs"
include "continuous/models_bjt.scs"
include "continuous/models_diodes.scs"
include "continuous/models_resistors.scs"
include "continuous/models_capacitors.scs"
include "corners/fs.scs"
include "corners/fs/specialized_cells.scs"
include "rescap/res_high__cap_low.scs"
include "rescap/res_high__cap_low__lin.scs"
endsection fs_hl

section fs_lh
parameters mc_mm_switch=0
parameters mc_pr_switch=0
parameters corner_factor=1
parameters process_mc_factor=1
parameters mismatch_factor=1
include "continuous/parameters_fet_fs.scs"
include "continuous/parameters_res_low.scs"
include "continuous/parameters_cap_high.scs"
include "continuous/models_global.scs"
include "continuous/models_fet.scs"
include "continuous/models_bjt.scs"
include "continuous/models_diodes.scs"
include "continuous/models_resistors.scs"
include "continuous/models_capacitors.scs"
include "corners/fs.scs"
include "corners/fs/specialized_cells.scs"
include "rescap/res_low__cap_high.scs"
include "rescap/res_low__cap_high__lin.scs"
endsection fs_lh

section fs_hh
parameters mc_mm_switch=0
parameters mc_pr_switch=0
parameters corner_factor=1
parameters process_mc_factor=1
parameters mismatch_factor=1
include "continuous/parameters_fet_fs.scs"
include "continuous/parameters_res_high.scs"
include "continuous/parameters_cap_high.scs"
include "continuous/models_global.scs"
include "continuous/models_fet.scs"
include "continuous/models_bjt.scs"
include "continuous/models_diodes.scs"
include "continuous/models_resistors.scs"
include "continuous/models_capacitors.scs"
include "corners/fs.scs"
include "corners/fs/specialized_cells.scs"
include "rescap/res_high__cap_high.scs"
include "rescap/res_high__cap_high__lin.scs"
endsection fs_hh

section ff_ll
parameters mc_mm_switch=0
parameters mc_pr_switch=0
parameters corner_factor=1
parameters process_mc_factor=1
parameters mismatch_factor=1
include "continuous/parameters_fet_ff.scs"
include "continuous/parameters_res_low.scs"
include "continuous/parameters_cap_low.scs"
include "continuous/models_global.scs"
include "continuous/models_fet.scs"
include "continuous/models_bjt.scs"
include "continuous/models_diodes.scs"
include "continuous/models_resistors.scs"
include "continuous/models_capacitors.scs"
include "corners/ff.scs"
include "corners/ff/specialized_cells.scs"
include "rescap/res_low__cap_low.scs"
include "rescap/res_low__cap_low__lin.scs"
endsection ff_ll

section ff_hl
parameters mc_mm_switch=0
parameters mc_pr_switch=0
parameters corner_factor=1
parameters process_mc_factor=1
parameters mismatch_factor=1
include "continuous/parameters_fet_ff.scs"
include "continuous/parameters_res_high.scs"
include "continuous/parameters_cap_low.scs"
include "continuous/models_global.scs"
include "continuous/models_fet.scs"
include "continuous/models_bjt.scs"
include "continuous/models_diodes.scs"
include "continuous/models_resistors.scs"
include "continuous/models_capacitors.scs"
include "corners/ff.scs"
include "corners/ff/specialized_cells.scs"
include "rescap/res_high__cap_low.scs"
include "rescap/res_high__cap_low__lin.scs"
endsection ff_hl

section ff_lh
parameters mc_mm_switch=0
parameters mc_pr_switch=0
parameters corner_factor=1
parameters process_mc_factor=1
parameters mismatch_factor=1
include "continuous/parameters_fet_ff.scs"
include "continuous/parameters_res_low.scs"
include "continuous/parameters_cap_high.scs"
include "continuous/models_global.scs"
include "continuous/models_fet.scs"
include "continuous/models_bjt.scs"
include "continuous/models_diodes.scs"
include "continuous/models_resistors.scs"
include "continuous/models_capacitors.scs"
include "corners/ff.scs"
include "corners/ff/specialized_cells.scs"
include "rescap/res_low__cap_high.scs"
include "rescap/res_low__cap_high__lin.scs"
endsection ff_lh

section ff_hh
parameters mc_mm_switch=0
parameters mc_pr_switch=0
parameters corner_factor=1
parameters process_mc_factor=1
parameters mismatch_factor=1
include "continuous/parameters_fet_ff.scs"
include "continuous/parameters_res_high.scs"
include "continuous/parameters_cap_high.scs"
include "continuous/models_global.scs"
include "continuous/models_fet.scs"
include "continuous/models_bjt.scs"
include "continuous/models_diodes.scs"
include "continuous/models_resistors.scs"
include "continuous/models_capacitors.scs"
include "corners/ff.scs"
include "corners/ff/specialized_cells.scs"
include "rescap/res_high__cap_high.scs"
include "rescap/res_high__cap_high__lin.scs"
endsection ff_hh

section tt_mm
parameters mc_mm_switch=1
parameters mc_pr_switch=0
parameters corner_factor=1
parameters process_mc_factor=1
parameters mismatch_factor=1
include "continuous/parameters_fet_tt.scs"
include "continuous/parameters_res_nom.scs"
include "continuous/parameters_cap_nom.scs"
include "continuous/models_global.scs"
include "continuous/models_fet.scs"
include "continuous/models_bjt.scs"
include "continuous/models_diodes.scs"
include "continuous/models_resistors.scs"
include "continuous/models_capacitors.scs"
include "corners/tt.scs"
include "corners/tt/specialized_cells.scs"
include "rescap/res_typical__cap_typical.scs"
include "rescap/res_typical__cap_typical__lin.scs"
endsection tt_mm

section sf_mm
parameters mc_mm_switch=1
parameters mc_pr_switch=0
parameters corner_factor=1
parameters process_mc_factor=1
parameters mismatch_factor=1
include "continuous/parameters_fet_sf.scs"
include "continuous/parameters_res_nom.scs"
include "continuous/parameters_cap_nom.scs"
include "continuous/models_global.scs"
include "continuous/models_fet.scs"
include "continuous/models_bjt.scs"
include "continuous/models_diodes.scs"
include "continuous/models_resistors.scs"
include "continuous/models_capacitors.scs"
include "corners/sf.scs"
include "corners/sf/specialized_cells.scs"
include "rescap/res_typical__cap_typical.scs"
include "rescap/res_typical__cap_typical__lin.scs"
endsection sf_mm

section ff_mm
parameters mc_mm_switch=1
parameters mc_pr_switch=0
parameters corner_factor=1
parameters process_mc_factor=1
parameters mismatch_factor=1
include "continuous/parameters_fet_ff.scs"
include "continuous/parameters_res_nom.scs"
include "continuous/parameters_cap_nom.scs"
include "continuous/models_global.scs"
include "continuous/models_fet.scs"
include "continuous/models_bjt.scs"
include "continuous/models_diodes.scs"
include "continuous/models_resistors.scs"
include "continuous/models_capacitors.scs"
include "corners/ff.scs"
include "corners/ff/specialized_cells.scs"
include "rescap/res_typical__cap_typical.scs"
include "rescap/res_typical__cap_typical__lin.scs"
endsection ff_mm

section ss_mm
parameters mc_mm_switch=1
parameters mc_pr_switch=0
parameters corner_factor=1
parameters process_mc_factor=1
parameters mismatch_factor=1
include "continuous/parameters_fet_ss.scs"
include "continuous/parameters_res_nom.scs"
include "continuous/parameters_cap_nom.scs"
include "continuous/models_global.scs"
include "continuous/models_fet.scs"
include "continuous/models_bjt.scs"
include "continuous/models_diodes.scs"
include "continuous/models_resistors.scs"
include "continuous/models_capacitors.scs"
include "corners/ss.scs"
include "corners/ss/specialized_cells.scs"
include "rescap/res_typical__cap_typical.scs"
include "rescap/res_typical__cap_typical__lin.scs"
endsection ss_mm

section fs_mm
parameters mc_mm_switch=1
parameters mc_pr_switch=0
parameters corner_factor=1
parameters process_mc_factor=1
parameters mismatch_factor=1
include "continuous/parameters_fet_fs.scs"
include "continuous/parameters_res_nom.scs"
include "continuous/parameters_cap_nom.scs"
include "continuous/models_global.scs"
include "continuous/models_fet.scs"
include "continuous/models_bjt.scs"
include "continuous/models_diodes.scs"
include "continuous/models_resistors.scs"
include "continuous/models_capacitors.scs"
include "corners/fs.scs"
include "corners/fs/specialized_cells.scs"
include "rescap/res_typical__cap_typical.scs"
include "rescap/res_typical__cap_typical__lin.scs"
endsection fs_mm

section ll_mm
parameters mc_mm_switch=1
parameters mc_pr_switch=0
parameters corner_factor=1
parameters process_mc_factor=1
parameters mismatch_factor=1
include "continuous/parameters_fet_tt.scs"
include "continuous/parameters_res_low.scs"
include "continuous/parameters_cap_low.scs"
include "continuous/models_global.scs"
include "continuous/models_fet.scs"
include "continuous/models_bjt.scs"
include "continuous/models_diodes.scs"
include "continuous/models_resistors.scs"
include "continuous/models_capacitors.scs"
include "corners/tt.scs"
include "corners/tt/specialized_cells.scs"
include "rescap/res_low__cap_low.scs"
include "rescap/res_low__cap_low__lin.scs"
endsection ll_mm

section hh_mm
parameters mc_mm_switch=1
parameters mc_pr_switch=0
parameters corner_factor=1
parameters process_mc_factor=1
parameters mismatch_factor=1
include "continuous/parameters_fet_tt.scs"
include "continuous/parameters_res_high.scs"
include "continuous/parameters_cap_high.scs"
include "continuous/models_global.scs"
include "continuous/models_fet.scs"
include "continuous/models_bjt.scs"
include "continuous/models_diodes.scs"
include "continuous/models_resistors.scs"
include "continuous/models_capacitors.scs"
include "corners/tt.scs"
include "corners/tt/specialized_cells.scs"
include "rescap/res_high__cap_high.scs"
include "rescap/res_high__cap_high__lin.scs"
endsection hh_mm

section hl_mm
parameters mc_mm_switch=1
parameters mc_pr_switch=0
parameters corner_factor=1
parameters process_mc_factor=1
parameters mismatch_factor=1
include "continuous/parameters_fet_tt.scs"
include "continuous/parameters_res_high.scs"
include "continuous/parameters_cap_low.scs"
include "continuous/models_global.scs"
include "continuous/models_fet.scs"
include "continuous/models_bjt.scs"
include "continuous/models_diodes.scs"
include "continuous/models_resistors.scs"
include "continuous/models_capacitors.scs"
include "corners/tt.scs"
include "corners/tt/specialized_cells.scs"
include "rescap/res_high__cap_low.scs"
include "rescap/res_high__cap_low__lin.scs"
endsection hl_mm

section lh_mm
parameters mc_mm_switch=1
parameters mc_pr_switch=0
parameters corner_factor=1
parameters process_mc_factor=1
parameters mismatch_factor=1
include "continuous/parameters_fet_tt.scs"
include "continuous/parameters_res_low.scs"
include "continuous/parameters_cap_high.scs"
include "continuous/models_global.scs"
include "continuous/models_fet.scs"
include "continuous/models_bjt.scs"
include "continuous/models_diodes.scs"
include "continuous/models_resistors.scs"
include "continuous/models_capacitors.scs"
include "corners/tt.scs"
include "corners/tt/specialized_cells.scs"
include "rescap/res_low__cap_high.scs"
include "rescap/res_low__cap_high__lin.scs"
endsection lh_mm

section ss_ll_mm
parameters mc_mm_switch=1
parameters mc_pr_switch=0
parameters corner_factor=1
parameters process_mc_factor=1
parameters mismatch_factor=1
include "continuous/parameters_fet_ss.scs"
include "continuous/parameters_res_low.scs"
include "continuous/parameters_cap_low.scs"
include "continuous/models_global.scs"
include "continuous/models_fet.scs"
include "continuous/models_bjt.scs"
include "continuous/models_diodes.scs"
include "continuous/models_resistors.scs"
include "continuous/models_capacitors.scs"
include "corners/ss.scs"
include "corners/ss/specialized_cells.scs"
include "rescap/res_low__cap_low.scs"
include "rescap/res_low__cap_low__lin.scs"
endsection ss_ll_mm

section ss_hl_mm
parameters mc_mm_switch=1
parameters mc_pr_switch=0
parameters corner_factor=1
parameters process_mc_factor=1
parameters mismatch_factor=1
include "continuous/parameters_fet_ss.scs"
include "continuous/parameters_res_high.scs"
include "continuous/parameters_cap_low.scs"
include "continuous/models_global.scs"
include "continuous/models_fet.scs"
include "continuous/models_bjt.scs"
include "continuous/models_diodes.scs"
include "continuous/models_resistors.scs"
include "continuous/models_capacitors.scs"
include "corners/ss.scs"
include "corners/ss/specialized_cells.scs"
include "rescap/res_high__cap_low.scs"
include "rescap/res_high__cap_low__lin.scs"
endsection ss_hl_mm

section ss_lh_mm
parameters mc_mm_switch=1
parameters mc_pr_switch=0
parameters corner_factor=1
parameters process_mc_factor=1
parameters mismatch_factor=1
include "continuous/parameters_fet_ss.scs"
include "continuous/parameters_res_low.scs"
include "continuous/parameters_cap_high.scs"
include "continuous/models_global.scs"
include "continuous/models_fet.scs"
include "continuous/models_bjt.scs"
include "continuous/models_diodes.scs"
include "continuous/models_resistors.scs"
include "continuous/models_capacitors.scs"
include "corners/ss.scs"
include "corners/ss/specialized_cells.scs"
include "rescap/res_low__cap_high.scs"
include "rescap/res_low__cap_high__lin.scs"
endsection ss_lh_mm

section ss_hh_mm
parameters mc_mm_switch=1
parameters mc_pr_switch=0
parameters corner_factor=1
parameters process_mc_factor=1
parameters mismatch_factor=1
include "continuous/parameters_fet_ss.scs"
include "continuous/parameters_res_high.scs"
include "continuous/parameters_cap_high.scs"
include "continuous/models_global.scs"
include "continuous/models_fet.scs"
include "continuous/models_bjt.scs"
include "continuous/models_diodes.scs"
include "continuous/models_resistors.scs"
include "continuous/models_capacitors.scs"
include "corners/ss.scs"
include "corners/ss/specialized_cells.scs"
include "rescap/res_high__cap_high.scs"
include "rescap/res_high__cap_high__lin.scs"
endsection ss_hh_mm

section sf_ll_mm
parameters mc_mm_switch=1
parameters mc_pr_switch=0
parameters corner_factor=1
parameters process_mc_factor=1
parameters mismatch_factor=1
include "continuous/parameters_fet_sf.scs"
include "continuous/parameters_res_low.scs"
include "continuous/parameters_cap_low.scs"
include "continuous/models_global.scs"
include "continuous/models_fet.scs"
include "continuous/models_bjt.scs"
include "continuous/models_diodes.scs"
include "continuous/models_resistors.scs"
include "continuous/models_capacitors.scs"
include "corners/sf.scs"
include "corners/sf/specialized_cells.scs"
include "rescap/res_low__cap_low.scs"
include "rescap/res_low__cap_low__lin.scs"
endsection sf_ll_mm

section sf_hl_mm
parameters mc_mm_switch=1
parameters mc_pr_switch=0
parameters corner_factor=1
parameters process_mc_factor=1
parameters mismatch_factor=1
include "continuous/parameters_fet_sf.scs"
include "continuous/parameters_res_high.scs"
include "continuous/parameters_cap_low.scs"
include "continuous/models_global.scs"
include "continuous/models_fet.scs"
include "continuous/models_bjt.scs"
include "continuous/models_diodes.scs"
include "continuous/models_resistors.scs"
include "continuous/models_capacitors.scs"
include "corners/sf.scs"
include "corners/sf/specialized_cells.scs"
include "rescap/res_high__cap_low.scs"
include "rescap/res_high__cap_low__lin.scs"
endsection sf_hl_mm

section sf_hh_mm
parameters mc_mm_switch=1
parameters mc_pr_switch=0
parameters corner_factor=1
parameters process_mc_factor=1
parameters mismatch_factor=1
include "continuous/parameters_fet_sf.scs"
include "continuous/parameters_res_high.scs"
include "continuous/parameters_cap_high.scs"
include "continuous/models_global.scs"
include "continuous/models_fet.scs"
include "continuous/models_bjt.scs"
include "continuous/models_diodes.scs"
include "continuous/models_resistors.scs"
include "continuous/models_capacitors.scs"
include "corners/sf.scs"
include "corners/sf/specialized_cells.scs"
include "rescap/res_high__cap_high.scs"
include "rescap/res_high__cap_high__lin.scs"
endsection sf_hh_mm

section fs_ll_mm
parameters mc_mm_switch=1
parameters mc_pr_switch=0
parameters corner_factor=1
parameters process_mc_factor=1
parameters mismatch_factor=1
include "continuous/parameters_fet_fs.scs"
include "continuous/parameters_res_low.scs"
include "continuous/parameters_cap_low.scs"
include "continuous/models_global.scs"
include "continuous/models_fet.scs"
include "continuous/models_bjt.scs"
include "continuous/models_diodes.scs"
include "continuous/models_resistors.scs"
include "continuous/models_capacitors.scs"
include "corners/fs.scs"
include "corners/fs/specialized_cells.scs"
include "rescap/res_low__cap_low.scs"
include "rescap/res_low__cap_low__lin.scs"
endsection fs_ll_mm

section fs_hl_mm
parameters mc_mm_switch=1
parameters mc_pr_switch=0
parameters corner_factor=1
parameters process_mc_factor=1
parameters mismatch_factor=1
include "continuous/parameters_fet_fs.scs"
include "continuous/parameters_res_high.scs"
include "continuous/parameters_cap_low.scs"
include "continuous/models_global.scs"
include "continuous/models_fet.scs"
include "continuous/models_bjt.scs"
include "continuous/models_diodes.scs"
include "continuous/models_resistors.scs"
include "continuous/models_capacitors.scs"
include "corners/fs.scs"
include "corners/fs/specialized_cells.scs"
include "rescap/res_high__cap_low.scs"
include "rescap/res_high__cap_low__lin.scs"
endsection fs_hl_mm

section fs_lh_mm
parameters mc_mm_switch=1
parameters mc_pr_switch=0
parameters corner_factor=1
parameters process_mc_factor=1
parameters mismatch_factor=1
include "continuous/parameters_fet_fs.scs"
include "continuous/parameters_res_low.scs"
include "continuous/parameters_cap_high.scs"
include "continuous/models_global.scs"
include "continuous/models_fet.scs"
include "continuous/models_bjt.scs"
include "continuous/models_diodes.scs"
include "continuous/models_resistors.scs"
include "continuous/models_capacitors.scs"
include "corners/fs.scs"
include "corners/fs/specialized_cells.scs"
include "rescap/res_low__cap_high.scs"
include "rescap/res_low__cap_high__lin.scs"
endsection fs_lh_mm

section fs_hh_mm
parameters mc_mm_switch=1
parameters mc_pr_switch=0
parameters corner_factor=1
parameters process_mc_factor=1
parameters mismatch_factor=1
include "continuous/parameters_fet_fs.scs"
include "continuous/parameters_res_high.scs"
include "continuous/parameters_cap_high.scs"
include "continuous/models_global.scs"
include "continuous/models_fet.scs"
include "continuous/models_bjt.scs"
include "continuous/models_diodes.scs"
include "continuous/models_resistors.scs"
include "continuous/models_capacitors.scs"
include "corners/fs.scs"
include "corners/fs/specialized_cells.scs"
include "rescap/res_high__cap_high.scs"
include "rescap/res_high__cap_high__lin.scs"
endsection fs_hh_mm

section ff_ll_mm
parameters mc_mm_switch=1
parameters mc_pr_switch=0
parameters corner_factor=1
parameters process_mc_factor=1
parameters mismatch_factor=1
include "continuous/parameters_fet_ff.scs"
include "continuous/parameters_res_low.scs"
include "continuous/parameters_cap_low.scs"
include "continuous/models_global.scs"
include "continuous/models_fet.scs"
include "continuous/models_bjt.scs"
include "continuous/models_diodes.scs"
include "continuous/models_resistors.scs"
include "continuous/models_capacitors.scs"
include "corners/ff.scs"
include "corners/ff/specialized_cells.scs"
include "rescap/res_low__cap_low.scs"
include "rescap/res_low__cap_low__lin.scs"
endsection ff_ll_mm

section ff_hl_mm
parameters mc_mm_switch=1
parameters mc_pr_switch=0
parameters corner_factor=1
parameters process_mc_factor=1
parameters mismatch_factor=1
include "continuous/parameters_fet_ff.scs"
include "continuous/parameters_res_high.scs"
include "continuous/parameters_cap_low.scs"
include "continuous/models_global.scs"
include "continuous/models_fet.scs"
include "continuous/models_bjt.scs"
include "continuous/models_diodes.scs"
include "continuous/models_resistors.scs"
include "continuous/models_capacitors.scs"
include "corners/ff.scs"
include "corners/ff/specialized_cells.scs"
include "rescap/res_high__cap_low.scs"
include "rescap/res_high__cap_low__lin.scs"
endsection ff_hl_mm

section ff_lh_mm
parameters mc_mm_switch=1
parameters mc_pr_switch=0
parameters corner_factor=1
parameters process_mc_factor=1
parameters mismatch_factor=1
include "continuous/parameters_fet_ff.scs"
include "continuous/parameters_res_low.scs"
include "continuous/parameters_cap_high.scs"
include "continuous/models_global.scs"
include "continuous/models_fet.scs"
include "continuous/models_bjt.scs"
include "continuous/models_diodes.scs"
include "continuous/models_resistors.scs"
include "continuous/models_capacitors.scs"
include "corners/ff.scs"
include "corners/ff/specialized_cells.scs"
include "rescap/res_low__cap_high.scs"
include "rescap/res_low__cap_high__lin.scs"
endsection ff_lh_mm

section ff_hh_mm
parameters mc_mm_switch=1
parameters mc_pr_switch=0
parameters corner_factor=1
parameters process_mc_factor=1
parameters mismatch_factor=1
include "continuous/parameters_fet_ff.scs"
include "continuous/parameters_res_high.scs"
include "continuous/parameters_cap_high.scs"
include "continuous/models_global.scs"
include "continuous/models_fet.scs"
include "continuous/models_bjt.scs"
include "continuous/models_diodes.scs"
include "continuous/models_resistors.scs"
include "continuous/models_capacitors.scs"
include "corners/ff.scs"
include "corners/ff/specialized_cells.scs"
include "rescap/res_high__cap_high.scs"
include "rescap/res_high__cap_high__lin.scs"
endsection ff_hh_mm

section mc
parameters mc_mm_switch=0
parameters mc_pr_switch=1
parameters corner_factor=1
parameters process_mc_factor=1
parameters mismatch_factor=1
include "continuous/parameters_fet_tt.scs"
include "continuous/parameters_res_nom.scs"
include "continuous/parameters_cap_nom.scs"
include "continuous/models_global.scs"
include "continuous/models_fet.scs"
include "continuous/models_bjt.scs"
include "continuous/models_diodes.scs"
include "continuous/models_resistors.scs"
include "continuous/models_capacitors.scs"
include "parameters/critical.scs"
include "parameters/montecarlo.scs"
endsection mc


endlibrary sky130.lib
