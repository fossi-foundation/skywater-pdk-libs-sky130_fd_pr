* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.include "models_fet/sky130_fd_pr__esd_nfet_05v0_nvt.spice"
.include "models_fet/sky130_fd_pr__esd_nfet_g5v0d10v5.spice"
.include "models_fet/sky130_fd_pr__esd_pfet_g5v0d10v5.spice"
.include "models_fet/sky130_fd_pr__nfet_01v8.spice"
.include "models_fet/sky130_fd_pr__nfet_01v8_esd.spice"
.include "models_fet/sky130_fd_pr__nfet_01v8_lvt.spice"
.include "models_fet/sky130_fd_pr__nfet_03v3_nvt.spice"
.include "models_fet/sky130_fd_pr__nfet_05v0_nvt.spice"
.include "models_fet/sky130_fd_pr__nfet_20v0.spice"
.include "models_fet/sky130_fd_pr__nfet_20v0_iso.spice"
.include "models_fet/sky130_fd_pr__nfet_20v0_nvt.spice"
.include "models_fet/sky130_fd_pr__nfet_20v0_zvt.spice"
.include "models_fet/sky130_fd_pr__nfet_g5v0d10v5.spice"
.include "models_fet/sky130_fd_pr__nfet_g5v0d16v0.spice"
.include "models_fet/sky130_fd_pr__nfet_g5v0d16v0_base.spice"
.include "models_fet/sky130_fd_pr__pfet_01v8.spice"
.include "models_fet/sky130_fd_pr__pfet_01v8_hvt.spice"
.include "models_fet/sky130_fd_pr__pfet_01v8_lvt.spice"
.include "models_fet/sky130_fd_pr__pfet_20v0.spice"
.include "models_fet/sky130_fd_pr__pfet_g5v0d10v5.spice"
.include "models_fet/sky130_fd_pr__pfet_g5v0d16v0.spice"
.include "models_fet/sky130_fd_pr__pfet_g5v0d16v0_base.spice"
