* SKY130 Spice File.
.param
+ tol_nfom=0
+ tol_pfom=0
+ tol_nw = 0.0
+ tol_poly = 0.0
+ tol_li = 0.0
+ tol_m1 = 0.0
+ tol_m2 = 0.0
+ tol_m3 = 0.0
+ tol_m4 = 0.0
+ tol_m5 = 0.0
+ tol_rdl = 0.0
.param
+ rcn=182
+ rcp=600
+ rdn=120
+ rdp=197
+ rdn_hv=114
+ rdp_hv=191
+ rp1=48.2
+ rnw=1700
+ rl1=12.2
+ rm1=0.125
+ rm2=0.125
+ rm3=0.047
+ rm4=0.047
+ rm5=0.0285
+ rrdl=0.005
+ rcp1=145.28
+ rcl1=9.3
+ rcvia=4.5
+ rcvia2=3.41
+ rcvia3=3.41
+ rcvia4=0.38
+ rcrdlcon=0.0058
+ rspwres=3816
* Interconnect Capacitance Parameters
.param
+ cp1f = 1.06e-04  cp1fsw = 8.64e-11
+ cl1f = 3.69e-05  cl1fsw = 8.30e-11
+ cl1d = 5.53e-05  cl1dsw = 8.23e-11
+ cl1p1 = 9.41e-05  cl1p1sw = 8.13e-11
+ cm1f = 2.58e-05  cm1fsw = 1.07e-10
+ cm1d = 3.36e-05  cm1dsw = 1.06e-10
+ cm1p1 = 4.48e-05  cm1p1sw = 1.06e-10
+ cm1l1 = 1.14e-04  cm1l1sw = 1.03e-10
+ cm2f = 1.75e-05  cm2fsw = 1.08e-10
+ cm2d = 2.08e-05  cm2dsw = 1.07e-10
+ cm2p1 = 2.47e-05  cm2p1sw = 1.07e-10
+ cm2l1 = 3.70e-05  cm2l1sw = 1.06e-10
+ cm2m1 = 1.28e-04  cm2m1sw = 1.03e-10
+ cm3f = 1.26e-05  cm3fsw = 1.08e-10
+ cm3d = 1.42e-05  cm3dsw = 1.09e-10
+ cm3p1 = 1.58e-05  cm3p1sw = 1.08e-10
+ cm3l1 = 2.02e-05  cm3l1sw = 1.08e-10
+ cm3m1 = 3.29e-05  cm3m1sw = 1.07e-10
+ cm3m2 = 8.22e-05  cm3m2sw = 1.05e-10
+ cm4f = 8.67e-06  cm4fsw = 1.09e-10
+ cm4d = 9.41e-06  cm4dsw = 1.09e-10
+ cm4p1 = 1.01e-05  cm4p1sw = 1.09e-10
+ cm4l1 = 1.17e-05  cm4l1sw = 1.09e-10
+ cm4m1 = 1.51e-05  cm4m1sw = 1.08e-10
+ cm4m2 = 2.09e-05  cm4m2sw = 1.08e-10
+ cm4m3 = 8.85e-05  cm4m3sw = 1.05e-10
+ cm5f = 6.48e-06  cm5fsw = 7.85e-11
+ cm5d = 6.88e-06  cm5dsw = 7.84e-11
+ cm5p1 = 7.26e-06  cm5p1sw = 7.82e-11
+ cm5l1 = 8.04e-06  cm5l1sw = 7.80e-11
+ cm5m1 = 9.50e-06  cm5m1sw = 7.77e-11
+ cm5m2 = 1.15e-05  cm5m2sw = 7.74e-11
+ cm5m3 = 1.99e-05  cm5m3sw = 7.76e-11
+ cm5m4 = 6.84e-05  cm5m4sw = 8.87e-11
+ crdlf = 2.57e-06  crdlfsw = 5.75e-11
+ crdld = 2.63e-06  crdldsw = 5.75e-11
+ crdlp1 = 2.68e-06  crdlp1sw = 5.74e-11
+ crdll1 = 2.78e-06  crdll1sw = 5.73e-11
+ crdlm1 = 2.93e-06  crdlm1sw = 5.71e-11
+ crdlm2 = 3.10e-06  crdlm2sw = 5.70e-11
+ crdlm3 = 3.50e-06  crdlm3sw = 5.68e-11
+ crdlm4 = 4.00e-06  crdlm4sw = 5.66e-11
+ crdlm5 = 5.44e-06  crdlm5sw = 5.68e-11
+ cl1p1f = 2.00e-04  cl1p1fsw = 8.32e-11
+ cm1p1f = 1.51e-04  cm1p1fsw = 8.45e-11
+ cm2p1f = 1.31e-04  cm2p1fsw = 8.53e-11
+ cm3p1f = 1.22e-04  cm3p1fsw = 8.58e-11
+ cm4p1f = 1.16e-04  cm4p1fsw = 8.61e-11
+ cm5p1f = 1.13e-04  cm5p1fsw = 8.61e-11
+ crdlp1f = 1.09e-04  crdlp1fsw = 8.63e-11
+ cm1l1f = 1.51e-04  cm1l1fsw = 7.90e-11
+ cm1l1d = 1.69e-04  cm1l1dsw = 7.81e-11
+ cm1l1p1 = 2.08e-04  cm1l1p1sw = 7.71e-11
+ cm2l1f = 7.40e-05  cm2l1fsw = 8.14e-11
+ cm2l1d = 9.23e-05  cm2l1dsw = 8.04e-11
+ cm2l1p1 = 1.31e-04  cm2l1p1sw = 7.94e-11
+ cm3l1f = 5.71e-05  cm3l1fsw = 8.21e-11
+ cm3l1d = 7.54e-05  cm3l1dsw = 8.13e-11
+ cm3l1p1 = 1.14e-04  cm3l1p1sw = 8.04e-11
+ cm4l1f = 4.86e-05  cm4l1fsw = 8.26e-11
+ cm4l1d = 6.70e-05  cm4l1dsw = 8.18e-11
+ cm4l1p1 = 1.06e-04  cm4l1p1sw = 8.08e-11
+ cm5l1f = 4.49e-05  cm5l1fsw = 8.28e-11
+ cm5l1d = 6.33e-05  cm5l1dsw = 8.20e-11
+ cm5l1p1 = 1.02e-04  cm5l1p1sw = 8.09e-11
+ crdll1f = 3.97e-05  crdll1fsw = 8.30e-11
+ crdll1d = 5.80e-05  crdll1dsw = 8.22e-11
+ crdll1p1 = 9.69e-05  crdll1p1sw = 8.12e-11
+ cm2m1f = 1.54e-04  cm2m1fsw = 1.02e-10
+ cm2m1d = 1.62e-04  cm2m1dsw = 1.02e-10
+ cm2m1p1 = 1.73e-04  cm2m1p1sw = 1.01e-10
+ cm2m1l1 = 2.42e-04  cm2m1l1sw = 9.89e-11
+ cm3m1f = 5.87e-05  cm3m1fsw = 1.05e-10
+ cm3m1d = 6.65e-05  cm3m1dsw = 1.04e-10
+ cm3m1p1 = 7.78e-05  cm3m1p1sw = 1.04e-10
+ cm3m1l1 = 1.47e-04  cm3m1l1sw = 1.02e-10
+ cm4m1f = 4.09e-05  cm4m1fsw = 1.07e-10
+ cm4m1d = 4.87e-05  cm4m1dsw = 1.06e-10
+ cm4m1p1 = 6.00e-05  cm4m1p1sw = 1.06e-10
+ cm4m1l1 = 1.29e-04  cm4m1l1sw = 1.03e-10
+ cm5m1f = 3.53e-05  cm5m1fsw = 1.07e-10
+ cm5m1d = 4.31e-05  cm5m1dsw = 1.06e-10
+ cm5m1p1 = 5.44e-05  cm5m1p1sw = 1.06e-10
+ cm5m1l1 = 1.23e-04  cm5m1l1sw = 1.04e-10
+ crdlm1f = 2.87e-05  crdlm1fsw = 1.07e-10
+ crdlm1d = 3.65e-05  crdlm1dsw = 1.07e-10
+ crdlm1p1 = 4.78e-05  crdlm1p1sw = 1.06e-10
+ crdlm1l1 = 1.17e-04  crdlm1l1sw = 1.03e-10
+ cm3m2f = 9.98e-05  cm3m2fsw = 1.03e-10
+ cm3m2d = 1.03e-04  cm3m2dsw = 1.03e-10
+ cm3m2p1 = 1.07e-04  cm3m2p1sw = 1.04e-10
+ cm3m2l1 = 1.19e-04  cm3m2l1sw = 1.02e-10
+ cm3m2m1 = 2.10e-04  cm3m2m1sw = 9.97e-11
+ cm4m2f = 3.84e-05  cm4m2fsw = 1.07e-10
+ cm4m2d = 4.17e-05  cm4m2dsw = 1.06e-10
+ cm4m2p1 = 4.56e-05  cm4m2p1sw = 1.06e-10
+ cm4m2l1 = 5.79e-05  cm4m2l1sw = 1.05e-10
+ cm4m2m1 = 1.49e-04  cm4m2m1sw = 1.03e-10
+ cm5m2f = 2.91e-05  cm5m2fsw = 1.07e-10
+ cm5m2d = 3.23e-05  cm5m2dsw = 1.07e-10
+ cm5m2p1 = 3.62e-05  cm5m2p1sw = 1.07e-10
+ cm5m2l1 = 4.85e-05  cm5m2l1sw = 1.05e-10
+ cm5m2m1 = 1.39e-04  cm5m2m1sw = 1.03e-10
+ crdlm2f = 2.06e-05  crdlm2fsw = 1.07e-10
+ crdlm2d = 2.39e-05  crdlm2dsw = 1.07e-10
+ crdlm2p1 = 2.78e-05  crdlm2p1sw = 1.07e-10
+ crdlm2l1 = 4.01e-05  crdlm2l1sw = 1.06e-10
+ crdlm2m1 = 1.31e-04  crdlm2m1sw = 1.03e-10
+ cm4m3f = 1.01e-04  cm4m3fsw = 1.03e-10
+ cm4m3d = 1.03e-04  cm4m3dsw = 1.03e-10
+ cm4m3p1 = 1.04e-04  cm4m3p1sw = 1.03e-10
+ cm4m3l1 = 1.09e-04  cm4m3l1sw = 1.03e-10
+ cm4m3m1 = 1.21e-04  cm4m3m1sw = 1.02e-10
+ cm4m3m2 = 1.71e-04  cm4m3m2sw = 9.99e-11
+ cm5m3f = 3.24e-05  cm5m3fsw = 1.06e-10
+ cm5m3d = 3.40e-05  cm5m3dsw = 1.06e-10
+ cm5m3p1 = 3.57e-05  cm5m3p1sw = 1.06e-10
+ cm5m3l1 = 4.00e-05  cm5m3l1sw = 1.05e-10
+ cm5m3m1 = 5.27e-05  cm5m3m1sw = 1.05e-10
+ cm5m3m2 = 1.02e-04  cm5m3m2sw = 1.03e-10
+ crdlm3f = 1.61e-05  crdlm3fsw = 1.08e-10
+ crdlm3d = 1.77e-05  crdlm3dsw = 1.08e-10
+ crdlm3p1 = 1.94e-05  crdlm3p1sw = 1.07e-10
+ crdlm3l1 = 2.37e-05  crdlm3l1sw = 1.07e-10
+ crdlm3m1 = 3.64e-05  crdlm3m1sw = 1.06e-10
+ crdlm3m2 = 8.57e-05  crdlm3m2sw = 1.05e-10
+ cm5m4f = 7.70e-05  cm5m4fsw = 1.04e-10
+ cm5m4d = 7.78e-05  cm5m4dsw = 1.04e-10
+ cm5m4p1 = 7.85e-05  cm5m4p1sw = 1.04e-10
+ cm5m4l1 = 8.01e-05  cm5m4l1sw = 1.04e-10
+ cm5m4m1 = 8.35e-05  cm5m4m1sw = 1.03e-10
+ cm5m4m2 = 8.92e-05  cm5m4m2sw = 1.03e-10
+ cm5m4m3 = 1.57e-04  cm5m4m3sw = 1.00e-10
+ crdlm4f = 1.27e-05  crdlm4fsw = 1.09e-10
+ crdlm4d = 1.34e-05  crdlm4dsw = 1.09e-10
+ crdlm4p1 = 1.41e-05  crdlm4p1sw = 1.09e-10
+ crdlm4l1 = 1.57e-05  crdlm4l1sw = 1.09e-10
+ crdlm4m1 = 1.91e-05  crdlm4m1sw = 1.08e-10
+ crdlm4m2 = 2.49e-05  crdlm4m2sw = 1.08e-10
+ crdlm4m3 = 9.25e-05  crdlm4m3sw = 1.05e-10
+ crdlm5f = 1.20e-05  crdlm5fsw = 7.60e-11
+ crdlm5d = 1.24e-05  crdlm5dsw = 7.59e-11
+ crdlm5p1 = 1.27e-05  crdlm5p1sw = 7.57e-11
+ crdlm5l1 = 1.35e-05  crdlm5l1sw = 7.55e-11
+ crdlm5m1 = 1.50e-05  crdlm5m1sw = 7.52e-11
+ crdlm5m2 = 1.70e-05  crdlm5m2sw = 7.49e-11
+ crdlm5m3 = 2.53e-05  crdlm5m3sw = 7.50e-11
+ crdlm5m4 = 7.39e-05  crdlm5m4sw = 8.61e-11
* P+ Poly Preres Parameters
.param
+ crpf_precision = 1.06e-04  ; Units: farad/meter^2
+ crpfsw_precision_1_1 = 5.04e-11 ; Units: farad/meter
+ crpfsw_precision_2_1 = 5.39e-11 ; Units: farad/meter
+ crpfsw_precision_4_1 = 5.83e-11 ; Units: farad/meter
+ crpfsw_precision_8_2 = 6.36e-11 ; Units: farad/meter
+ crpfsw_precision_16_2 = 6.97e-11 ; Units: farad/meter
.include "sky130_fd_pr__model__res.model.spice"
