* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

******************************************************************
******************************************************************
*  *****************************************************
*  04/14/2021 Usman Suriono
*      Why     : New scalable sky130_fd_pr__nfet_01v8 native 3V model
*      What    : Converted from discrete ntvnative model
*      What    : Converted from discrete nshort model
*                Replaced rsh from 1 to calculated rsh from the original model.
*                PDK netlist nrd/nrs = ratio of distance the middle of the contact to Gate.
*
*  *****************************************************
*
*  Nmos Native 3V Model
*  -----------------------------------------------------

.subckt  sky130_fd_pr__nfet_03v3_nvt  d g s b  mult=1
+ 
.param  l = 1 w = 1 nf = 1 ad = 0 as = 0 pd = 0 ps = 0 nrd = {0.14/w} nrs = {0.14/w} sa = 0 sb = 0 sd = 0
+ swx_nrds = {89.1*nf/w+443.5}
+ swx_vth = {sw_vth0_sky130_fd_pr__nfet_01v8_nat+sw_mm_vth0_sky130_fd_pr__nfet_01v8_nat*mismatch_factor*MC_MM_SWITCH*AGAUSS(0,1.0,1)/sqrt(l*w*mult)+sw_vth0_sky130_fd_pr__nfet_01v8_nat_mc}

Msky130_fd_pr__nfet_03v3_nvt  d g s b ntvnative_model l = {l} w = {w} ad = {ad} as = {as} pd = {pd} ps = {ps} nrd = {nrd} nrs = {nrs} sa = {sa} sb = {sb} sd = {sd} nf = {nf}
* + deltox = 0.3*(sw_tox_hv_corner - sw_tox_hv_nom) + sw_tox_hv_mc + sw_mm_tox_hv * mismatch_factor*MC_MM_SWITCH*AGAUSS(0,1.0,1)/sqrt(l*w*mult)
* + mulu0  = sw_u0_sky130_fd_pr__nfet_01v8_nat**(1.3*(0.22*10/w+0.78))
* + mulvsat= 0.85
+ delvto = {-0.0387+1.37*swx_vth*(0.026*10/w+0.974)+0.0058/w}




.model ntvnative_model.1 nmos
+ level = 54 lmin = 6E-7 lmax = 9.079999999999999E-7 wmin = 4E-6
+ wmax = 1.01E-4 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 1.16E-8
+ toxm = 1.16E-8 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 9.999999999999999E22 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0.01855708
+ wint = {1E-8+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {5E-8-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = 0 dwb = 0 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = 0.0713243 k1 = 0.33502
+ k2 = 5.7767E-3 k3 = -0.5 k3b = 0
+ w0 = 0 lpe0 = -1E-10 lpeb = 0
+ vbm = -3 dvtp0 = 0 dvtp1 = 0
+ dvt0 = 1E-10 dvt1 = 0.536 dvt2 = -0.05
+ dvt0w = 0 dvt1w = 5E6 dvt2w = -0.032
+ vfbsdoff = 0 u0 = 0.0898544 ua = 4.203204E-9
+ ub = 2.98748E-18 uc = 1.3541E-10 ud = 0
+ up = 0 lp = 1 eu = 1.67
+ vsat = 1.139932E5 a0 = 3.1139121E-4 ags = 1.4554757E-4
+ b0 = 0 b1 = 0 keta = -0.016684
+ a1 = 0 a2 = 0.6218093 rdsw = 0
+ rdswmin = 0 rdw = 0 rdwmin = 0
+ rsw = 0 rswmin = 0 prwb = 0
+ prwg = 0 wr = 1 voff = -0.098774
+ voffl = -2.9752837E-11 minv = 0 nfactor = 0.30842
+ eta0 = 0 etab = 0 dsub = 0.071143
+ cit = -3.3686011E-37 cdsc = 0 cdscb = -1E-4
+ cdscd = 1.5E-5 pclm = 2.8944111 pdiblc1 = 0.87012255
+ pdiblc2 = 0.032974 pdiblcb = -0.05 drout = 0.27268
+ pscbe1 = 4.24E9 pscbe2 = 1E-8 pvag = 5.2718232
+ delta = 0.01 fprout = 10.125 pdits = 5.666761E-16
+ pditsl = 0 pditsd = 0 lambda = 0
+ vtl = 0 lc = 5E-9 xn = 3
+ alpha0 = 8.3952E-7 alpha1 = 0.33 beta0 = 23
+ aigbacc = 0.43 bigbacc = 0.054 cigbacc = 0.075
+ nigbacc = 1 aigbinv = 0.35 bigbinv = 0.03
+ cigbinv = 6E-3 eigbinv = 1.1 nigbinv = 3
+ aigc = 0.43 bigc = 0.054 cigc = 0.075
+ aigsd = 0.43 bigsd = 0.054 cigsd = 0.075
+ dlcig = 0 nigc = 1 poxedge = 1
+ pigcd = 1 ntox = 1 toxref = 1.16E-8
+ agidl = 0 bgidl = 2.3E9 cgidl = 0.8
+ egidl = 0.5 noia = 2.5E41 noib = 0
+ noic = 0 em = 4.1E7 af = 1
+ ef = 1 kf = 0 lintnoi = 0
+ tnoia = 6.4E6 tnoib = 7.2E6 ntnoi = 1
+ rnoia = 0.89 rnoib = 0.38 xpart = 0
+ cgso = {2.517561582E-10/sw_func_tox_hv_ratio} cgdo = {2.517561582E-10/sw_func_tox_hv_ratio} cgbo = {0/sw_func_tox_hv_ratio}
+ ckappas = 0.6 cf = 0 clc = 1E-7
+ cle = 0.6 dlc = 4.9452E-8 dwc = 0
+ vfbcv = -1 noff = 4 voffcv = -0.14208
+ acde = 0.4 moin = 15 cgsl = {3.85585E-11/sw_func_tox_hv_ratio}
+ cgdl = {3.85585E-11/sw_func_tox_hv_ratio} ijthsrev = 0.1 ijthsfwd = 0.1
+ xjbvs = 1 bvs = 12.69 jss = 4.2966E-4
+ jsws = 8.040000000000001E-10 cjs = {8.310E-04*sw_func_nsd_pw_cj} mjs = 0.28329
+ mjsws = 0.057926 cjsws = {8.88731424E-11*sw_func_nsd_pw_cj} cjswgs = {3.736446E-11*sw_func_nsd_pw_cj}
+ mjswgs = 0.33 pbs = 0.66345 pbsws = 1
+ pbswgs = 0.2442 xrcrg1 = 12 xrcrg2 = 1
+ rbpb = 50 rbpd = 50 rbps = 50
+ rbdb = 50 rbsb = 50 gbmin = 1E-12
+ tnom = 30 ute = -1.613 kt1 = -0.29818
+ kt1l = 0 kt2 = -0.02 ua1 = 1E-9
+ ub1 = -8.411E-18 uc1 = -2.5133E-10 at = 3.726E4
+ prt = 0 njs = 1.5764 xtis = 0
+ tpb = 1.9685E-3 tpbsw = 1E-3 tpbswg = 0
+ tcj = 8.3E-4 tcjsw = 0 tcjswg = 0
+ tvoff = 0 tvfbsdoff = 0 saref = 1.95E-6
+ sbref = 1.94E-6 wlod = 0 ku0 = -3E-8
+ kvsat = 0.3 kvth0 = -2E-9 tku0 = 0
+ llodku0 = 0 wlodku0 = 1 llodvth = 0
+ wlodvth = 1 lku0 = 0 wku0 = 5E-7
+ pku0 = 0 lkvth0 = 0 wkvth0 = 0
+ pkvth0 = 0 stk2 = 0 lodk2 = 1
+ steta0 = 0 lodeta0 = 1

.model ntvnative_model.2 nmos
+ level = 54 lmin = 5E-7 lmax = 6E-7 wmin = 4E-6
+ wmax = 1.01E-4 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 1.16E-8
+ toxm = 1.16E-8 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 9.999999999999999E22 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0.01855708
+ wint = {1E-8+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {5E-8-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = 0 dwb = 0 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = 0.501080966666667 lvth0 = -2.57854E-7
+ wvth0 = 9.713333333333337E-8 pvth0 = -5.828000000000002E-14 k1 = 0.66012
+ lk1 = -1.9506E-7 k2 = 0.029621366666667 lk2 = -1.43068E-8
+ wk2 = -4.528666666666667E-8 pk2 = 2.7172E-14 k3 = -0.5
+ k3b = 0 w0 = 0 lpe0 = -1E-10
+ lpeb = 0 vbm = -3 dvtp0 = 0
+ dvtp1 = 0 dvt0 = 1E-10 dvt1 = 0.536
+ dvt2 = -0.05 dvt0w = 0 dvt1w = 5E6
+ dvt2w = -0.032 vfbsdoff = 0 u0 = 0.07427035
+ lu0 = 9.350430000000007E-9 wu0 = 1.038590000000002E-7 pu0 = -6.231540000000009E-14
+ ua = -1.426761E-9 lua = 3.377979E-15 wua = 4.835999999999991E-15
+ pua = -2.901599999999994E-21 ub = 1.770416333333334E-17 lub = -8.830010000000002E-24
+ wub = 6.409666666666668E-24 pub = -3.845800000000001E-30 uc = 1.3541E-10
+ ud = 0 up = 0 lp = 1
+ eu = 1.67 vsat = 1.276985333333333E5 lvsat = -8.223199999999986E-3
+ wvsat = -0.048033333333333 pvsat = 2.882000000000001E-8 a0 = 3.1139121E-4
+ ags = 1.4554757E-4 b0 = 0 b1 = 0
+ keta = -0.135433 lketa = 7.124940000000003E-8 a1 = 0
+ a2 = 0.6218093 rdsw = 0 rdswmin = 0
+ rdw = 0 rdwmin = 0 rsw = 0
+ rswmin = 0 prwb = 0 prwg = 0
+ wr = 1 voff = -0.283605666666667 lvoff = 1.10899E-7
+ wvoff = -7.413333333333348E-8 pvoff = 4.448000000000009E-14 voffl = -2.9752837E-11
+ minv = 0 nfactor = -1.335146666666667 lnfactor = 9.8614E-7
+ wnfactor = -7.233333333333352E-7 pnfactor = 4.340000000000012E-13 eta0 = -0.08669
+ leta0 = 5.201400000000001E-8 etab = 0 dsub = -2.537442000000001
+ ldsub = 1.565151000000001E-6 cit = -3.3686011E-37 cdsc = 0
+ cdscb = -1E-4 cdscd = 1.5E-5 pclm = 2.8944111
+ pdiblc1 = 0.87012255 pdiblc2 = 0.032974 pdiblcb = -0.05
+ drout = 0.27268 pscbe1 = 4.24E9 pscbe2 = 1E-8
+ pvag = 5.2718232 delta = 0.01 fprout = 10.125
+ pdits = 5.666761E-16 pditsl = 0 pditsd = 0
+ lambda = 0 vtl = 0 lc = 5E-9
+ xn = 3 alpha0 = 2.407320000000001E-6 lalpha0 = -9.406800000000006E-13
+ walpha0 = -4.872000000000003E-12 palpha0 = 2.923200000000002E-18 alpha1 = 1.980000000000001
+ lalpha1 = -9.900000000000003E-7 beta0 = 30.870000000000005 lbeta0 = -4.722000000000002E-6
+ wbeta0 = -1.940000000000003E-5 pbeta0 = 1.164000000000002E-11 aigbacc = 0.43
+ bigbacc = 0.054 cigbacc = 0.075 nigbacc = 1
+ aigbinv = 0.35 bigbinv = 0.03 cigbinv = 6E-3
+ eigbinv = 1.1 nigbinv = 3 aigc = 0.43
+ bigc = 0.054 cigc = 0.075 aigsd = 0.43
+ bigsd = 0.054 cigsd = 0.075 dlcig = 0
+ nigc = 1 poxedge = 1 pigcd = 1
+ ntox = 1 toxref = 1.16E-8 agidl = 0
+ bgidl = 2.3E9 cgidl = 0.8 egidl = 0.5
+ noia = 2.5E41 noib = 0 noic = 0
+ em = 4.1E7 af = 1 ef = 1
+ kf = 0 lintnoi = 0 tnoia = 6.4E6
+ tnoib = 7.2E6 ntnoi = 1 rnoia = 0.89
+ rnoib = 0.38 xpart = 0 cgso = {2.517561582E-10/sw_func_tox_hv_ratio}
+ cgdo = {2.517561582E-10/sw_func_tox_hv_ratio} cgbo = {0/sw_func_tox_hv_ratio} ckappas = 0.6
+ cf = 0 clc = 1E-7 cle = 0.6
+ dlc = 4.9452E-8 dwc = 0 vfbcv = -1
+ noff = 4 voffcv = -0.14208 acde = 0.4
+ moin = 15 cgsl = {3.85585E-11/sw_func_tox_hv_ratio} cgdl = {3.85585E-11/sw_func_tox_hv_ratio}
+ ijthsrev = 0.1 ijthsfwd = 0.1 xjbvs = 1
+ bvs = 12.69 jss = 4.2966E-4 jsws = 8.040000000000001E-10
+ cjs = {8.310E-04*sw_func_nsd_pw_cj} mjs = 0.28329 mjsws = 0.057926
+ cjsws = {8.88731424E-11*sw_func_nsd_pw_cj} cjswgs = {3.736446E-11*sw_func_nsd_pw_cj} mjswgs = 0.33
+ pbs = 0.66345 pbsws = 1 pbswgs = 0.2442
+ xrcrg1 = 12 xrcrg2 = 1 rbpb = 50
+ rbpd = 50 rbps = 50 rbdb = 50
+ rbsb = 50 gbmin = 1E-12 tnom = 30
+ ute = -1.098 lute = -3.09E-7 kt1 = -0.09488
+ lkt1 = -1.2198E-7 kt1l = 0 kt2 = -0.186666666666667
+ lkt2 = 1E-7 wkt2 = 6.666666666666669E-7 pkt2 = -4.000000000000001E-13
+ ua1 = 1E-9 ub1 = 5.387333333333346E-18 lub1 = -8.279000000000006E-24
+ wub1 = 3.146666666666664E-23 pub1 = -1.887999999999998E-29 uc1 = 7.342533333333335E-10
+ luc1 = -5.913500000000001E-16 wuc1 = -3.942333333333335E-15 puc1 = 2.365400000000001E-21
+ at = 2.105999999999999E4 lat = 9.720000000000003E-3 prt = 0
+ njs = 1.5764 xtis = 0 tpb = 1.9685E-3
+ tpbsw = 1E-3 tpbswg = 0 tcj = 8.3E-4
+ tcjsw = 0 tcjswg = 0 tvoff = 0
+ tvfbsdoff = 0 saref = 1.95E-6 sbref = 1.94E-6
+ wlod = 0 ku0 = -3E-8 kvsat = 0.3
+ kvth0 = -2E-9 tku0 = 0 llodku0 = 0
+ wlodku0 = 1 llodvth = 0 wlodvth = 1
+ lku0 = 0 wku0 = 5E-7 pku0 = 0
+ lkvth0 = 0 wkvth0 = 0 pkvth0 = 0
+ stk2 = 0 lodk2 = 1 steta0 = 0
+ lodeta0 = 1

.model ntvnative_model.3 nmos
+ level = 54 lmin = 6E-7 lmax = 9.079999999999999E-7 wmin = 1E-6
+ wmax = 4E-6 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 1.16E-8
+ toxm = 1.16E-8 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 9.999999999999999E22 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0.01855708
+ wint = {1E-8+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {5E-8-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = 0 dwb = 0 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = 0.0713243 k1 = 0.33502
+ k2 = 5.7767E-3 k3 = -0.5 k3b = 0
+ w0 = 0 lpe0 = -1E-10 lpeb = 0
+ vbm = -3 dvtp0 = 0 dvtp1 = 0
+ dvt0 = 1E-10 dvt1 = 0.536 dvt2 = -0.05
+ dvt0w = 0 dvt1w = 5E6 dvt2w = -0.032
+ vfbsdoff = 0 u0 = 0.0898544 ua = 4.203204E-9
+ ub = 2.98748E-18 uc = 1.3541E-10 ud = 0
+ up = 0 lp = 1 eu = 1.67
+ vsat = 1.139932E5 a0 = 3.1139121E-4 ags = 1.4554757E-4
+ b0 = 0 b1 = 0 keta = -0.016684
+ a1 = 0 a2 = 0.6218093 rdsw = 0
+ rdswmin = 0 rdw = 0 rdwmin = 0
+ rsw = 0 rswmin = 0 prwb = 0
+ prwg = 0 wr = 1 voff = -0.098774
+ voffl = -2.9752837E-11 minv = 0 nfactor = 0.30842
+ eta0 = 0 etab = 0 dsub = 0.071143
+ cit = -3.3686011E-37 cdsc = 0 cdscb = -1E-4
+ cdscd = 1.5E-5 pclm = 2.8944111 pdiblc1 = 0.87012255
+ pdiblc2 = 0.032974 pdiblcb = -0.05 drout = 0.27268
+ pscbe1 = 4.24E9 pscbe2 = 1E-8 pvag = 5.2718232
+ delta = 0.01 fprout = 10.125 pdits = 5.666761E-16
+ pditsl = 0 pditsd = 0 lambda = 0
+ vtl = 0 lc = 5E-9 xn = 3
+ alpha0 = 8.3952E-7 alpha1 = 0.33 beta0 = 23
+ aigbacc = 0.43 bigbacc = 0.054 cigbacc = 0.075
+ nigbacc = 1 aigbinv = 0.35 bigbinv = 0.03
+ cigbinv = 6E-3 eigbinv = 1.1 nigbinv = 3
+ aigc = 0.43 bigc = 0.054 cigc = 0.075
+ aigsd = 0.43 bigsd = 0.054 cigsd = 0.075
+ dlcig = 0 nigc = 1 poxedge = 1
+ pigcd = 1 ntox = 1 toxref = 1.16E-8
+ agidl = 0 bgidl = 2.3E9 cgidl = 0.8
+ egidl = 0.5 noia = 2.5E41 noib = 0
+ noic = 0 em = 4.1E7 af = 1
+ ef = 1 kf = 0 lintnoi = 0
+ tnoia = 6.4E6 tnoib = 7.2E6 ntnoi = 1
+ rnoia = 0.89 rnoib = 0.38 xpart = 0
+ cgso = {2.517561582E-10/sw_func_tox_hv_ratio} cgdo = {2.517561582E-10/sw_func_tox_hv_ratio} cgbo = {0/sw_func_tox_hv_ratio}
+ ckappas = 0.6 cf = 0 clc = 1E-7
+ cle = 0.6 dlc = 4.9452E-8 dwc = 0
+ vfbcv = -1 noff = 4 voffcv = -0.14208
+ acde = 0.4 moin = 15 cgsl = {3.85585E-11/sw_func_tox_hv_ratio}
+ cgdl = {3.85585E-11/sw_func_tox_hv_ratio} ijthsrev = 0.1 ijthsfwd = 0.1
+ xjbvs = 1 bvs = 12.69 jss = 4.2966E-4
+ jsws = 8.040000000000001E-10 cjs = {8.310E-04*sw_func_nsd_pw_cj} mjs = 0.28329
+ mjsws = 0.057926 cjsws = {8.88731424E-11*sw_func_nsd_pw_cj} cjswgs = {3.736446E-11*sw_func_nsd_pw_cj}
+ mjswgs = 0.33 pbs = 0.66345 pbsws = 1
+ pbswgs = 0.2442 xrcrg1 = 12 xrcrg2 = 1
+ rbpb = 50 rbpd = 50 rbps = 50
+ rbdb = 50 rbsb = 50 gbmin = 1E-12
+ tnom = 30 ute = -1.613 kt1 = -0.29818
+ kt1l = 0 kt2 = -0.02 ua1 = 1E-9
+ ub1 = -8.411E-18 uc1 = -2.5133E-10 at = 3.726E4
+ prt = 0 njs = 1.5764 xtis = 0
+ tpb = 1.9685E-3 tpbsw = 1E-3 tpbswg = 0
+ tcj = 8.3E-4 tcjsw = 0 tcjswg = 0
+ tvoff = 0 tvfbsdoff = 0 saref = 1.95E-6
+ sbref = 1.94E-6 wlod = 0 ku0 = -3E-8
+ kvsat = 0.3 kvth0 = -2E-9 tku0 = 0
+ llodku0 = 0 wlodku0 = 1 llodvth = 0
+ wlodvth = 1 lku0 = 0 wku0 = 5E-7
+ pku0 = 0 lkvth0 = 0 wkvth0 = 0
+ pkvth0 = 0 stk2 = 0 lodk2 = 1
+ steta0 = 0 lodeta0 = 1

.model ntvnative_model.4 nmos
+ level = 54 lmin = 5E-7 lmax = 6E-7 wmin = 1E-6
+ wmax = 4E-6 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 1.16E-8
+ toxm = 1.16E-8 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 9.999999999999999E22 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0.01855708
+ wint = {1E-8+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {5E-8-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = 0 dwb = 0 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = 0.5310743 lvth0 = -2.7585E-7
+ wvth0 = -2.284E-8 pvth0 = 1.3704E-14 k1 = 0.66012
+ lk1 = -1.9506E-7 k2 = 0.028970033333333 lk2 = -1.3916E-8
+ wk2 = -4.268133333333334E-8 pk2 = 2.56088E-14 k3 = -0.5
+ k3b = 0 w0 = 0 lpe0 = -1E-10
+ lpeb = 0 vbm = -3 dvtp0 = 0
+ dvtp1 = 0 dvt0 = 1E-10 dvt1 = 0.536
+ dvt2 = -0.05 dvt0w = 0 dvt1w = 5E6
+ dvt2w = -0.032 vfbsdoff = 0 u0 = 0.098487333333333
+ lu0 = -5.17976000000002E-9 wu0 = 6.991066666666622E-9 pu0 = -4.194639999999973E-15
+ ua = -5.277443333333358E-10 lua = 2.838569000000002E-15 wua = 1.23993333333334E-15
+ pua = -7.439600000000038E-22 ub = 2.003641333333334E-17 lub = -1.022936E-23
+ wub = -2.919333333333335E-24 pub = 1.751600000000001E-30 uc = 1.3541E-10
+ ud = 0 up = 0 lp = 1
+ eu = 1.67 vsat = 1.235442E5 lvsat = -5.730599999999979E-3
+ wvsat = -0.031416 pvsat = 1.884959999999998E-8 a0 = 3.1139121E-4
+ ags = 1.4554757E-4 b0 = 0 b1 = 0
+ keta = -0.115436 lketa = 5.925120000000002E-8 wketa = -7.998800000000003E-8
+ pketa = 4.799280000000001E-14 a1 = 0 a2 = 0.6218093
+ rdsw = 0 rdswmin = 0 rdw = 0
+ rdwmin = 0 rsw = 0 rswmin = 0
+ prwb = 0 prwg = 0 wr = 1
+ voff = -0.314790666666667 lvoff = 1.2961E-7 wvoff = 5.060666666666668E-8
+ pvoff = -3.036400000000001E-14 voffl = -2.9752837E-11 minv = 0
+ nfactor = -1.572146666666667 lnfactor = 1.12834E-6 wnfactor = 2.246666666666672E-7
+ pnfactor = -1.348000000000003E-13 eta0 = -0.112697 leta0 = 6.761820000000001E-8
+ weta0 = 1.04028E-7 peta0 = -6.241680000000001E-14 etab = 1.666666666666667E-10
+ letab = -1E-16 wetab = -6.666666666666668E-16 petab = 4.000000000000001E-22
+ dsub = -2.537442000000001 ldsub = 1.565151000000001E-6 cit = -3.3686011E-37
+ cdsc = 0 cdscb = -1E-4 cdscd = 1.5E-5
+ pclm = 2.8944111 pdiblc1 = 0.87012255 pdiblc2 = 0.032974
+ pdiblcb = -0.05 drout = 0.27268 pscbe1 = 4.24E9
+ pscbe2 = 1E-8 pvag = 5.2718232 delta = 0.01
+ fprout = 10.125 pdits = 5.666761E-16 pditsl = 0
+ pditsd = 0 lambda = 0 vtl = 0
+ lc = 5E-9 xn = 3 alpha0 = 7.229200000000002E-7
+ lalpha0 = 6.995999999999994E-14 walpha0 = 1.8656E-12 palpha0 = -1.11936E-18
+ alpha1 = 2.030000000000001 lalpha1 = -1.02E-6 walpha1 = -1.999999999999998E-7
+ palpha1 = 1.199999999999999E-13 beta0 = 23.393333333333324 lbeta0 = -2.359999999999967E-7
+ wbeta0 = 1.050666666666667E-5 pbeta0 = -6.304000000000004E-12 aigbacc = 0.43
+ bigbacc = 0.054 cigbacc = 0.075 nigbacc = 1
+ aigbinv = 0.35 bigbinv = 0.03 cigbinv = 6E-3
+ eigbinv = 1.1 nigbinv = 3 aigc = 0.43
+ bigc = 0.054 cigc = 0.075 aigsd = 0.43
+ bigsd = 0.054 cigsd = 0.075 dlcig = 0
+ nigc = 1 poxedge = 1 pigcd = 1
+ ntox = 1 toxref = 1.16E-8 agidl = 0
+ bgidl = 2.3E9 cgidl = 0.8 egidl = 0.5
+ noia = 2.5E41 noib = 0 noic = 0
+ em = 4.1E7 af = 1 ef = 1
+ kf = 0 lintnoi = 0 tnoia = 6.4E6
+ tnoib = 7.2E6 ntnoi = 1 rnoia = 0.89
+ rnoib = 0.38 xpart = 0 cgso = {2.517561582E-10/sw_func_tox_hv_ratio}
+ cgdo = {2.517561582E-10/sw_func_tox_hv_ratio} cgbo = {0/sw_func_tox_hv_ratio} ckappas = 0.6
+ cf = 0 clc = 1E-7 cle = 0.6
+ dlc = 4.9452E-8 dwc = 0 vfbcv = -1
+ noff = 4 voffcv = -0.14208 acde = 0.4
+ moin = 15 cgsl = {3.85585E-11/sw_func_tox_hv_ratio} cgdl = {3.85585E-11/sw_func_tox_hv_ratio}
+ ijthsrev = 0.1 ijthsfwd = 0.1 xjbvs = 1
+ bvs = 12.69 jss = 4.2966E-4 jsws = 8.040000000000001E-10
+ cjs = {8.310E-04*sw_func_nsd_pw_cj} mjs = 0.28329 mjsws = 0.057926
+ cjsws = {8.88731424E-11*sw_func_nsd_pw_cj} cjswgs = {3.736446E-11*sw_func_nsd_pw_cj} mjswgs = 0.33
+ pbs = 0.66345 pbsws = 1 pbswgs = 0.2442
+ xrcrg1 = 12 xrcrg2 = 1 rbpb = 50
+ rbpd = 50 rbps = 50 rbdb = 50
+ rbsb = 50 gbmin = 1E-12 tnom = 30
+ ute = -1.098 lute = -3.09E-7 kt1 = -0.09488
+ lkt1 = -1.2198E-7 kt1l = 0 kt2 = -0.02
+ ua1 = 1E-9 ub1 = 1.325400000000001E-17 lub1 = -1.2999E-23
+ uc1 = -2.5133E-10 at = 2.105999999999999E4 lat = 9.720000000000003E-3
+ prt = 0 njs = 1.5764 xtis = 0
+ tpb = 1.9685E-3 tpbsw = 1E-3 tpbswg = 0
+ tcj = 8.3E-4 tcjsw = 0 tcjswg = 0
+ tvoff = 0 tvfbsdoff = 0 saref = 1.95E-6
+ sbref = 1.94E-6 wlod = 0 ku0 = -3E-8
+ kvsat = 0.3 kvth0 = -2E-9 tku0 = 0
+ llodku0 = 0 wlodku0 = 1 llodvth = 0
+ wlodvth = 1 lku0 = 0 wku0 = 5E-7
+ pku0 = 0 lkvth0 = 0 wkvth0 = 0
+ pkvth0 = 0 stk2 = 0 lodk2 = 1
+ steta0 = 0 lodeta0 = 1

.model ntvnative_model.5 nmos
+ level = 54 lmin = 6E-7 lmax = 9.079999999999999E-7 wmin = 7E-7
+ wmax = 1E-6 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 1.16E-8
+ toxm = 1.16E-8 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 9.999999999999999E22 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0.01855708
+ wint = {1E-8+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {5E-8-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = 0 dwb = 0 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = 0.079979566666667 wvth0 = -8.655266666666637E-9
+ k1 = 0.33502 k2 = -5.302999999999974E-4 wk2 = 6.306999999999998E-9
+ k3 = -0.5 k3b = 0 w0 = 0
+ lpe0 = -1E-10 lpeb = 0 vbm = -3
+ dvtp0 = 0 dvtp1 = 0 dvt0 = 1E-10
+ dvt1 = 0.536 dvt2 = -0.05 dvt0w = 0
+ dvt1w = 5E6 dvt2w = -0.032 vfbsdoff = 0
+ u0 = 0.090725666666667 wu0 = -8.712666666666571E-10 ua = 4.200525E-9
+ ub = 3.325813333333333E-18 wub = -3.383333333333333E-25 uc = 1.3541E-10
+ ud = 0 up = 0 lp = 1
+ eu = 1.67 vsat = 1.110814333333333E5 wvsat = 2.911766666666687E-3
+ a0 = 3.1139121E-4 ags = 1.4554757E-4 b0 = 0
+ b1 = 0 keta = -0.0667746 wketa = 5.009059999999999E-8
+ a1 = 0 a2 = 0.6218093 rdsw = 0
+ rdswmin = 0 rdw = 0 rdwmin = 0
+ rsw = 0 rswmin = 0 prwb = 0
+ prwg = 0 wr = 1 voff = -0.098774
+ voffl = -2.9752837E-11 minv = 0 nfactor = 0.243576666666667
+ wnfactor = 6.484333333333328E-8 eta0 = 0 etab = 0
+ dsub = 0.071143 cit = -3.3686011E-37 cdsc = 0
+ cdscb = -1E-4 cdscd = 1.5E-5 pclm = 2.8944111
+ pdiblc1 = 0.87012255 pdiblc2 = 0.032974 pdiblcb = -0.05
+ drout = 0.27268 pscbe1 = 4.24E9 pscbe2 = 1E-8
+ pvag = 5.2718232 delta = 0.01 fprout = 10.125
+ pdits = 5.666761E-16 pditsl = 0 pditsd = 0
+ lambda = 0 vtl = 0 lc = 5E-9
+ xn = 3 alpha0 = 1.982199999999999E-6 walpha0 = -1.14268E-12
+ alpha1 = 0.283333333333333 walpha1 = 4.666666666666657E-8 beta0 = 26.308666666666664
+ wbeta0 = -3.308666666666664E-6 aigbacc = 0.43 bigbacc = 0.054
+ cigbacc = 0.075 nigbacc = 1 aigbinv = 0.35
+ bigbinv = 0.03 cigbinv = 6E-3 eigbinv = 1.1
+ nigbinv = 3 aigc = 0.43 bigc = 0.054
+ cigc = 0.075 aigsd = 0.43 bigsd = 0.054
+ cigsd = 0.075 dlcig = 0 nigc = 1
+ poxedge = 1 pigcd = 1 ntox = 1
+ toxref = 1.16E-8 agidl = 0 bgidl = 2.3E9
+ cgidl = 0.8 egidl = 0.5 noia = 2.5E41
+ noib = 0 noic = 0 em = 4.1E7
+ af = 1 ef = 1 kf = 0
+ lintnoi = 0 tnoia = 6.4E6 tnoib = 7.2E6
+ ntnoi = 1 rnoia = 0.89 rnoib = 0.38
+ xpart = 0 cgso = {2.517561582E-10/sw_func_tox_hv_ratio} cgdo = {2.517561582E-10/sw_func_tox_hv_ratio}
+ cgbo = {0/sw_func_tox_hv_ratio} ckappas = 0.6 cf = 0
+ clc = 1E-7 cle = 0.6 dlc = 4.9452E-8
+ dwc = 0 vfbcv = -1 noff = 4
+ voffcv = -0.14208 acde = 0.4 moin = 15
+ cgsl = {3.85585E-11/sw_func_tox_hv_ratio} cgdl = {3.85585E-11/sw_func_tox_hv_ratio} ijthsrev = 0.1
+ ijthsfwd = 0.1 xjbvs = 1 bvs = 12.69
+ jss = 4.2966E-4 jsws = 8.040000000000001E-10 cjs = {8.310E-04*sw_func_nsd_pw_cj}
+ mjs = 0.28329 mjsws = 0.057926 cjsws = {8.88731424E-11*sw_func_nsd_pw_cj}
+ cjswgs = {3.736446E-11*sw_func_nsd_pw_cj} mjswgs = 0.33 pbs = 0.66345
+ pbsws = 1 pbswgs = 0.2442 xrcrg1 = 12
+ xrcrg2 = 1 rbpb = 50 rbpd = 50
+ rbps = 50 rbdb = 50 rbsb = 50
+ gbmin = 1E-12 tnom = 30 ute = -1.4527
+ wute = -1.603E-7 kt1 = -0.28236 wkt1 = -1.582000000000002E-8
+ kt1l = 0 kt2 = -0.02 ua1 = 1E-9
+ ub1 = -4.842633333333333E-18 wub1 = -3.568366666666666E-24 uc1 = -2.5133E-10
+ at = 4.293E4 wat = -5.669999999999999E-3 prt = 0
+ njs = 1.5764 xtis = 0 tpb = 1.9685E-3
+ tpbsw = 1E-3 tpbswg = 0 tcj = 8.3E-4
+ tcjsw = 0 tcjswg = 0 tvoff = 0
+ tvfbsdoff = 0 saref = 1.95E-6 sbref = 1.94E-6
+ wlod = 0 ku0 = -3E-8 kvsat = 0.3
+ kvth0 = -2E-9 tku0 = 0 llodku0 = 0
+ wlodku0 = 1 llodvth = 0 wlodvth = 1
+ lku0 = 0 wku0 = 5E-7 pku0 = 0
+ lkvth0 = 0 wkvth0 = 0 pkvth0 = 0
+ stk2 = 0 lodk2 = 1 steta0 = 0
+ lodeta0 = 1

.model ntvnative_model.6 nmos
+ level = 54 lmin = 5E-7 lmax = 6E-7 wmin = 7E-7
+ wmax = 1E-6 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 1.16E-8
+ toxm = 1.16E-8 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 9.999999999999999E22 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0.01855708
+ wint = {1E-8+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {5E-8-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = 0 dwb = 0 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = 0.448594066666667 lvth0 = -2.211687E-7
+ wvth0 = 5.964023333333348E-8 pvth0 = -4.097730000000006E-14 k1 = 0.78612
+ lk1 = -2.706599999999998E-7 wk1 = -1.259999999999997E-7 pk1 = 7.559999999999984E-14
+ k2 = -0.0347218 lk2 = 2.05149E-8 wk2 = 2.10105E-8
+ pk2 = -8.8221E-15 k3 = -0.5 k3b = 0
+ w0 = 0 lpe0 = -1E-10 lpeb = 0
+ vbm = -3 dvtp0 = 0 dvtp1 = 0
+ dvt0 = 1E-10 dvt1 = 0.536 dvt2 = -0.05
+ dvt0w = 0 dvt1w = 5E6 dvt2w = -0.032
+ vfbsdoff = 0 u0 = 0.062575166666667 lu0 = 1.689030000000006E-8
+ wu0 = 4.290323333333345E-8 pu0 = -2.626470000000006E-14 ua = -3.93034166666665E-9
+ lua = 4.88387799999999E-15 wua = 4.642530666666652E-15 pua = -2.789268999999992E-21
+ ub = 2.129477333333334E-17 lub = -1.0781376E-23 wub = -4.177693333333336E-24
+ pub = 2.303616000000001E-30 uc = -6.228883333333333E-10 luc = 4.549789999999999E-16
+ wuc = 7.582983333333335E-16 puc = -4.54979E-22 ud = 0
+ up = 0 lp = 1 eu = 1.67
+ vsat = 9.50812666666666E4 lvsat = 9.600100000000025E-3 wvsat = -2.953066666666614E-3
+ pvsat = 3.51889999999998E-9 a0 = 3.1139121E-4 ags = 1.4554757E-4
+ b0 = 0 b1 = 0 keta = -0.4959676
+ lketa = 2.575158E-7 wketa = 3.005436E-7 pketa = -1.502718E-13
+ a1 = 0 a2 = 0.6218093 rdsw = 0
+ rdswmin = 0 rdw = 0 rdwmin = 0
+ rsw = 0 rswmin = 0 prwb = 0
+ prwg = 0 wr = 1 voff = -0.160957333333333
+ lvoff = 3.731000000000009E-8 wvoff = -1.032266666666666E-7 pvoff = 6.193599999999996E-14
+ voffl = -2.9752837E-11 minv = 0 nfactor = -1.127539999999999
+ lnfactor = 8.226699999999997E-7 wnfactor = -2.199400000000006E-7 pnfactor = 1.708700000000003E-13
+ eta0 = -0.0264693 leta0 = 1.588158E-8 weta0 = 1.78003E-8
+ peta0 = -1.068018E-14 etab = -5.000000000000001E-10 letab = 3.000000000000001E-16
+ dsub = -2.537442000000001 ldsub = 1.565151000000001E-6 cit = -3.3686011E-37
+ cdsc = 0 cdscb = -1E-4 cdscd = 1.5E-5
+ pclm = 2.8944111 pdiblc1 = 0.87012255 pdiblc2 = 0.032974
+ pdiblcb = -0.05 drout = 0.27268 pscbe1 = 4.24E9
+ pscbe2 = 1E-8 pvag = 5.2718232 delta = 0.01
+ fprout = 10.125 pdits = 5.666761E-16 pditsl = 0
+ pditsd = 0 lambda = 0 vtl = 0
+ lc = 5E-9 xn = 3 alpha0 = 8.383516666666669E-6
+ lalpha0 = -3.84079E-12 walpha0 = -5.794996666666667E-12 palpha0 = 2.79139E-18
+ alpha1 = 2.950000000000001 lalpha1 = -1.6E-6 walpha1 = -1.120000000000001E-6
+ palpha1 = 7.000000000000002E-13 beta0 = 48.38533333333332 lbeta0 = -1.324599999999999E-5
+ wbeta0 = -1.448533333333332E-5 pbeta0 = 6.705999999999989E-12 aigbacc = 0.43
+ bigbacc = 0.054 cigbacc = 0.075 nigbacc = 1
+ aigbinv = 0.35 bigbinv = 0.03 cigbinv = 6E-3
+ eigbinv = 1.1 nigbinv = 3 aigc = 0.43
+ bigc = 0.054 cigc = 0.075 aigsd = 0.43
+ bigsd = 0.054 cigsd = 0.075 dlcig = 0
+ nigc = 1 poxedge = 1 pigcd = 1
+ ntox = 1 toxref = 1.16E-8 agidl = 0
+ bgidl = 2.3E9 cgidl = 0.8 egidl = 0.5
+ noia = 2.5E41 noib = 0 noic = 0
+ em = 4.1E7 af = 1 ef = 1
+ kf = 0 lintnoi = 0 tnoia = 6.4E6
+ tnoib = 7.2E6 ntnoi = 1 rnoia = 0.89
+ rnoib = 0.38 xpart = 0 cgso = {2.517561582E-10/sw_func_tox_hv_ratio}
+ cgdo = {2.517561582E-10/sw_func_tox_hv_ratio} cgbo = {0/sw_func_tox_hv_ratio} ckappas = 0.6
+ cf = 0 clc = 1E-7 cle = 0.6
+ dlc = 4.9452E-8 dwc = 0 vfbcv = -1
+ noff = 4 voffcv = -0.14208 acde = 0.4
+ moin = 15 cgsl = {3.85585E-11/sw_func_tox_hv_ratio} cgdl = {3.85585E-11/sw_func_tox_hv_ratio}
+ ijthsrev = 0.1 ijthsfwd = 0.1 xjbvs = 1
+ bvs = 12.69 jss = 4.2966E-4 jsws = 8.040000000000001E-10
+ cjs = {8.310E-04*sw_func_nsd_pw_cj} mjs = 0.28329 mjsws = 0.057926
+ cjsws = {8.88731424E-11*sw_func_nsd_pw_cj} cjswgs = {3.736446E-11*sw_func_nsd_pw_cj} mjswgs = 0.33
+ pbs = 0.66345 pbsws = 1 pbswgs = 0.2442
+ xrcrg1 = 12 xrcrg2 = 1 rbpb = 50
+ rbpd = 50 rbps = 50 rbdb = 50
+ rbsb = 50 gbmin = 1E-12 tnom = 30
+ ute = 1.065466666666667 lute = -1.5109E-6 wute = -2.163466666666666E-6
+ pute = 1.2019E-12 kt1 = -0.07906 lkt1 = -1.2198E-7
+ wkt1 = -1.582000000000002E-8 kt1l = 0 kt2 = -0.02
+ ua1 = 1E-9 ub1 = 4.656419999999999E-17 lub1 = -3.084409999999999E-23
+ wub1 = -3.331019999999999E-23 pub1 = 1.784509999999999E-29 uc1 = -2.5133E-10
+ at = 5.507999999999999E4 lat = -7.289999999999999E-3 wat = -0.03402
+ pat = 1.701E-8 prt = 0 njs = 1.5764
+ xtis = 0 tpb = 1.9685E-3 tpbsw = 1E-3
+ tpbswg = 0 tcj = 8.3E-4 tcjsw = 0
+ tcjswg = 0 tvoff = 0 tvfbsdoff = 0
+ saref = 1.95E-6 sbref = 1.94E-6 wlod = 0
+ ku0 = -3E-8 kvsat = 0.3 kvth0 = -2E-9
+ tku0 = 0 llodku0 = 0 wlodku0 = 1
+ llodvth = 0 wlodvth = 1 lku0 = 0
+ wku0 = 5E-7 pku0 = 0 lkvth0 = 0
+ wkvth0 = 0 pkvth0 = 0 stk2 = 0
+ lodk2 = 1 steta0 = 0 lodeta0 = 1

.model ntvnative_model.7 nmos
+ level = 54 lmin = 6E-7 lmax = 9.079999999999999E-7 wmin = 4.2E-7
+ wmax = 7E-7 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 1.16E-8
+ toxm = 1.16E-8 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 9.999999999999999E22 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0.01855708
+ wint = {1E-8+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {5E-8-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = 0 dwb = 0 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = -0.12221325 lvth0 = 1.212804E-7
+ wvth0 = 1.32879705E-7 pvth0 = -8.489627999999998E-14 k1 = -0.046145
+ lk1 = 2.245319999999999E-7 wk1 = 2.668154999999999E-7 pk1 = -1.571723999999999E-13
+ k2 = 6.020750000000001E-3 lk2 = -2.336400000000001E-9 wk2 = 1.721265E-9
+ pk2 = 1.63548E-15 k3 = -0.5 k3b = 0
+ w0 = 0 lpe0 = -1E-10 lpeb = 0
+ vbm = -3 dvtp0 = 0 dvtp1 = 0
+ dvt0 = 1E-10 dvt1 = 0.536 dvt2 = -0.05
+ dvt0w = 0 dvt1w = 5E6 dvt2w = -0.032
+ vfbsdoff = 0 u0 = 0.1428645 lu0 = -3.299399999999998E-8
+ wu0 = -3.736844999999997E-8 pu0 = 2.309579999999998E-14 ua = 9.396800999999994E-9
+ lua = -2.800555199999997E-15 wua = -3.637393199999997E-15 pua = 1.960388639999998E-21
+ ub = 4.4244955E-18 lub = -1.1849724E-24 wub = -1.10741085E-24
+ pub = 8.2948068E-31 uc = 1.79915E-10 luc = 3.914279999999998E-17
+ wuc = -3.115350000000003E-17 puc = -2.739995999999998E-23 ud = 0
+ up = 0 lp = 1 eu = 1.67
+ vsat = 1.4699775E5 lvsat = -0.02419812 wvsat = -0.022229655
+ pvsat = 1.693868399999999E-8 a0 = 3.1139121E-4 ags = 1.4554757E-4
+ b0 = 0 b1 = 0 keta = 0.02019395
+ lketa = -6.588360000000001E-9 wketa = -1.0787385E-8 pketa = 4.611852E-15
+ a1 = 0 a2 = 0.6218093 rdsw = 0
+ rdswmin = 0 rdw = 0 rdwmin = 0
+ rsw = 0 rswmin = 0 prwb = 0
+ prwg = 0 wr = 1 voff = -0.098774
+ voffl = -2.9752837E-11 minv = 0 nfactor = 2.439824999999999
+ lnfactor = -1.31238E-6 wnfactor = -1.4725305E-6 pnfactor = 9.186659999999999E-13
+ eta0 = 9.362699999999997E-4 leta0 = -7.490159999999998E-10 weta0 = -6.553889999999998E-10
+ peta0 = 5.243111999999999E-16 etab = 4.499999999999998E-10 letab = -3.599999999999999E-16
+ wetab = -3.149999999999999E-16 petab = 2.52E-22 dsub = 2.4188695
+ ldsub = -1.8781812E-6 wdsub = -1.64340855E-6 pdsub = 1.31472684E-12
+ cit = -3.3686011E-37 cdsc = 0 cdscb = -1E-4
+ cdscd = 1.5E-5 pclm = 2.8944111 pdiblc1 = 0.87012255
+ pdiblc2 = 0.032974 pdiblcb = -0.05 drout = 0.27268
+ pscbe1 = 4.24E9 pscbe2 = 1E-8 pvag = 5.2718232
+ delta = 0.01 fprout = 10.125 pdits = 5.666761E-16
+ pditsl = 0 pditsd = 0 lambda = 0
+ vtl = 0 lc = 5E-9 xn = 3
+ alpha0 = -1.851599999999999E-6 lalpha0 = 1.153296E-12 walpha0 = 1.54098E-12
+ palpha0 = -8.073071999999998E-19 alpha1 = 0.335 lalpha1 = 3.239999999999999E-7
+ walpha1 = 1.049999999999989E-8 palpha1 = -2.268E-13 beta0 = 16.854000000000006
+ lbeta0 = 3.293999999999996E-6 wbeta0 = 3.309599999999996E-6 pbeta0 = -2.305799999999997E-12
+ aigbacc = 0.43 bigbacc = 0.054 cigbacc = 0.075
+ nigbacc = 1 aigbinv = 0.35 bigbinv = 0.03
+ cigbinv = 6E-3 eigbinv = 1.1 nigbinv = 3
+ aigc = 0.43 bigc = 0.054 cigc = 0.075
+ aigsd = 0.43 bigsd = 0.054 cigsd = 0.075
+ dlcig = 0 nigc = 1 poxedge = 1
+ pigcd = 1 ntox = 1 toxref = 1.16E-8
+ agidl = 0 bgidl = 2.3E9 cgidl = 0.8
+ egidl = 0.5 noia = 2.5E41 noib = 0
+ noic = 0 em = 4.1E7 af = 1
+ ef = 1 kf = 0 lintnoi = 0
+ tnoia = 6.4E6 tnoib = 7.2E6 ntnoi = 1
+ rnoia = 0.89 rnoib = 0.38 xpart = 0
+ cgso = {2.517561582E-10/sw_func_tox_hv_ratio} cgdo = {2.517561582E-10/sw_func_tox_hv_ratio} cgbo = {0/sw_func_tox_hv_ratio}
+ ckappas = 0.6 cf = 0 clc = 1E-7
+ cle = 0.6 dlc = 4.9452E-8 dwc = 0
+ vfbcv = -1 noff = 4 voffcv = -0.14208
+ acde = 0.4 moin = 15 cgsl = {3.85585E-11/sw_func_tox_hv_ratio}
+ cgdl = {3.85585E-11/sw_func_tox_hv_ratio} ijthsrev = 0.1 ijthsfwd = 0.1
+ xjbvs = 1 bvs = 12.69 jss = 4.2966E-4
+ jsws = 8.040000000000001E-10 cjs = {8.310E-04*sw_func_nsd_pw_cj} mjs = 0.28329
+ mjsws = 0.057926 cjsws = {8.88731424E-11*sw_func_nsd_pw_cj} cjswgs = {3.736446E-11*sw_func_nsd_pw_cj}
+ mjswgs = 0.33 pbs = 0.66345 pbsws = 1
+ pbswgs = 0.2442 xrcrg1 = 12 xrcrg2 = 1
+ rbpb = 50 rbpd = 50 rbps = 50
+ rbdb = 50 rbsb = 50 gbmin = 1E-12
+ tnom = 30 ute = -1.47605 lute = -2.469599999999999E-7
+ wute = -1.439549999999999E-7 pute = 1.728719999999999E-13 kt1 = -0.45742
+ lkt1 = 1.219679999999999E-7 wkt1 = 1.067219999999999E-7 pkt1 = -8.53775999999999E-14
+ kt1l = 0 kt2 = -0.02 ua1 = 1E-9
+ ub1 = -2.255649999999999E-17 lub1 = 6.422759999999997E-24 wub1 = 8.831339999999997E-24
+ pub1 = -4.495931999999998E-30 uc1 = -9.7517E-10 luc1 = 4.34304E-16
+ wuc1 = 5.06688E-16 puc1 = -3.040128E-22 at = 9.9225E4
+ lat = -0.04374 wat = -0.0450765 pat = 3.0618E-8
+ prt = 0 njs = 1.5764 xtis = 0
+ tpb = 1.9685E-3 tpbsw = 1E-3 tpbswg = 0
+ tcj = 8.3E-4 tcjsw = 0 tcjswg = 0
+ tvoff = 0 tvfbsdoff = 0 saref = 2.34E-6
+ sbref = 2.34E-6 wlod = 0 ku0 = -3E-8
+ kvsat = 0.3 kvth0 = -2E-9 tku0 = 0
+ llodku0 = 0 wlodku0 = 1 llodvth = 0
+ wlodvth = 1 lku0 = 0 wku0 = 5E-7
+ pku0 = 0 lkvth0 = 0 wkvth0 = 0
+ pkvth0 = 0 stk2 = 0 lodk2 = 1
+ steta0 = 0 lodeta0 = 1

.model ntvnative_model.8 nmos
+ level = 54 lmin = 5E-7 lmax = 6E-7 wmin = 4.2E-7
+ wmax = 7E-7 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 1.16E-8
+ toxm = 1.16E-8 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 9.999999999999999E22 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0.01855708
+ wint = {1E-8+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {5E-8-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = 0 dwb = 0 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = 0.490247 lvth0 = -2.461957500000001E-7
+ wvth0 = 3.048317999999996E-8 pvth0 = -2.345836499999998E-14 k1 = 0.7329
+ lk1 = -2.428949999999998E-7 wk1 = -8.874599999999978E-8 pk1 = 5.616449999999988E-14
+ k2 = -0.051172 lk2 = 3.197925000000001E-8 wk2 = 3.252564000000001E-8
+ pk2 = -1.6847145E-14 k3 = -0.5 k3b = 0
+ w0 = 0 lpe0 = -1E-10 lpeb = 0
+ vbm = -3 dvtp0 = 0 dvtp1 = 0
+ dvt0 = 1E-10 dvt1 = 0.536 dvt2 = -0.05
+ dvt0w = 0 dvt1w = 5E6 dvt2w = -0.032
+ vfbsdoff = 0 u0 = 0.11335125 lu0 = -1.528605000000008E-8
+ wu0 = 7.359974999999917E-9 pu0 = -3.741254999999957E-15 ua = 3.064501499999998E-9
+ lua = 9.988245000000013E-16 wua = -2.538595500000004E-16 pua = -6.97315499999999E-23
+ ub = 1.3541274E-17 lub = -6.6550395E-24 wub = 1.249756200000002E-24
+ pub = -5.848195500000011E-31 uc = 7.491855000000002E-10 luc = -3.024195E-16
+ wuc = -2.0215335E-16 puc = 7.519994999999999E-23 ud = 0
+ up = 0 lp = 1 eu = 1.67
+ vsat = 7.419954999999996E4 lvsat = 0.0194808 wvsat = 0.011664135
+ pvsat = -3.397590000000019E-9 a0 = 3.1139121E-4 ags = 1.4554757E-4
+ b0 = 0 b1 = 0 keta = 0.0457451
+ lketa = -2.191905000000002E-8 wketa = -7.865529000000002E-8 pketa = 4.533259500000001E-14
+ a1 = 0 a2 = 0.6218093 rdsw = 0
+ rdswmin = 0 rdw = 0 rdwmin = 0
+ rsw = 0 rswmin = 0 prwb = 0
+ prwg = 0 wr = 1 voff = -0.2820015
+ lvoff = 1.099365E-7 wvoff = -1.849575E-8 pvoff = 1.109745E-14
+ voffl = -2.9752837E-11 minv = 0 nfactor = -1.919850000000001
+ lnfactor = 1.303425E-6 wnfactor = 3.346770000000002E-7 pnfactor = -1.656585000000001E-13
+ eta0 = -2.91284E-3 leta0 = 1.56045E-9 weta0 = 1.310778E-9
+ peta0 = -6.553890000000002E-16 etab = -1.4E-9 letab = 7.500000000000003E-16
+ wetab = 6.300000000000001E-16 petab = -3.150000000000001E-22 dsub = -7.232895000000004
+ ldsub = 3.912877500000002E-6 wdsub = 3.286817100000002E-6 pdsub = -1.643408550000001E-12
+ cit = -3.3686011E-37 cdsc = 0 cdscb = -1E-4
+ cdscd = 1.5E-5 pclm = 2.8944111 pdiblc1 = 0.87012255
+ pdiblc2 = 0.032974 pdiblcb = -0.05 drout = 0.27268
+ pscbe1 = 4.24E9 pscbe2 = 1E-8 pvag = 5.2718232
+ delta = 0.01 fprout = 10.125 pdits = 5.666761E-16
+ pditsl = 0 pditsd = 0 lambda = 0
+ vtl = 0 lc = 5E-9 xn = 3
+ alpha0 = -4.937900000000003E-7 lalpha0 = 3.386100000000002E-13 walpha0 = 4.191180000000002E-13
+ palpha0 = -1.341900000000001E-19 alpha1 = 3.374999999999999 lalpha1 = -1.5E-6
+ walpha1 = -1.4175E-6 palpha1 = 6.300000000000001E-13 beta0 = 38.369
+ lbeta0 = -9.615000000000002E-6 wbeta0 = -7.473899999999996E-6 pbeta0 = 4.164299999999998E-12
+ aigbacc = 0.43 bigbacc = 0.054 cigbacc = 0.075
+ nigbacc = 1 aigbinv = 0.35 bigbinv = 0.03
+ cigbinv = 6E-3 eigbinv = 1.1 nigbinv = 3
+ aigc = 0.43 bigc = 0.054 cigc = 0.075
+ aigsd = 0.43 bigsd = 0.054 cigsd = 0.075
+ dlcig = 0 nigc = 1 poxedge = 1
+ pigcd = 1 ntox = 1 toxref = 1.16E-8
+ agidl = 0 bgidl = 2.3E9 cgidl = 0.8
+ egidl = 0.5 noia = 2.5E41 noib = 0
+ noic = 0 em = 4.1E7 af = 1
+ ef = 1 kf = 0 lintnoi = 0
+ tnoia = 6.4E6 tnoib = 7.2E6 ntnoi = 1
+ rnoia = 0.89 rnoib = 0.38 xpart = 0
+ cgso = {2.517561582E-10/sw_func_tox_hv_ratio} cgdo = {2.517561582E-10/sw_func_tox_hv_ratio} cgbo = {0/sw_func_tox_hv_ratio}
+ ckappas = 0.6 cf = 0 clc = 1E-7
+ cle = 0.6 dlc = 4.9452E-8 dwc = 0
+ vfbcv = -1 noff = 4 voffcv = -0.14208
+ acde = 0.4 moin = 15 cgsl = {3.85585E-11/sw_func_tox_hv_ratio}
+ cgdl = {3.85585E-11/sw_func_tox_hv_ratio} ijthsrev = 0.1 ijthsfwd = 0.1
+ xjbvs = 1 bvs = 12.69 jss = 4.2966E-4
+ jsws = 8.040000000000001E-10 cjs = {8.310E-04*sw_func_nsd_pw_cj} mjs = 0.28329
+ mjsws = 0.057926 cjsws = {8.88731424E-11*sw_func_nsd_pw_cj} cjswgs = {3.736446E-11*sw_func_nsd_pw_cj}
+ mjswgs = 0.33 pbs = 0.66345 pbsws = 1
+ pbswgs = 0.2442 xrcrg1 = 12 xrcrg2 = 1
+ rbpb = 50 rbpd = 50 rbps = 50
+ rbdb = 50 rbsb = 50 gbmin = 1E-12
+ tnom = 30 ute = -2.7464 lute = 5.1525E-7
+ wute = 5.0484E-7 pute = -2.16405E-13 kt1 = 0.152485
+ lkt1 = -2.439749999999998E-7 wkt1 = -1.779014999999998E-7 pkt1 = 8.539649999999992E-14
+ kt1l = 0 kt2 = -0.02 ua1 = 1E-9
+ ub1 = 4.70910000000001E-18 lub1 = -9.936600000000007E-24 wub1 = -4.011630000000004E-24
+ pub1 = 3.209850000000003E-30 uc1 = 7.288450000000003E-10 luc1 = -5.881050000000001E-16
+ wuc1 = -6.861225000000001E-16 puc1 = 4.116735000000001E-22 at = -4.455000000000002E4
+ lat = 0.042525 wat = 0.035721 pat = -1.78605E-8
+ prt = 0 njs = 1.5764 xtis = 0
+ tpb = 1.9685E-3 tpbsw = 1E-3 tpbswg = 0
+ tcj = 8.3E-4 tcjsw = 0 tcjswg = 0
+ tvoff = 0 tvfbsdoff = 0 saref = 1.95E-6
+ sbref = 1.94E-6 wlod = 0 ku0 = -3E-8
+ kvsat = 0.3 kvth0 = -2E-9 tku0 = 0
+ llodku0 = 0 wlodku0 = 1 llodvth = 0
+ wlodvth = 1 lku0 = 0 wku0 = 5E-7
+ pku0 = 0 lkvth0 = 0 wkvth0 = 0
+ pkvth0 = 0 stk2 = 0 lodk2 = 1
+ steta0 = 0 lodeta0 = 1

.ends sky130_fd_pr__nfet_03v3_nvt
