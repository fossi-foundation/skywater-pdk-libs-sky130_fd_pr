* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

******************************************************************
******************************************************************
*  *****************************************************
*  04/14/2021 Usman Suriono
*      Why     : New scalable sky130_fd_pr__pfet_01v8 low VT model
*      What    : Converted from discrete plowvt models
*                Replaced rsh from 1 to calculated rsh from the original model.
*                PDK netlist nrd/nrs = ratio of distance the middle of the contact to Gate.
*
*  *****************************************************
*
*  Pmos Low VT Model
*  -----------------------------------------------------

.subckt  sky130_fd_pr__pfet_01v8_lvt  d g s b  mult=1
+ 
.param  l = 1 w = 1 nf = 1 ad = 0 as = 0 pd = 0 ps = 0 nrd = {0.14/w} nrs = {0.14/w} sa = 0 sb = 0 sd = 0
+ swx_nrds = {361*nf/w+1489}

Msky130_fd_pr__pfet_01v8_lvt  d g s b plowvt_model l = {l} w = {w} ad = {ad} as = {as} pd = {pd} ps = {ps} nrd = {nrd} nrs = {nrs} sa = {sa} sb = {sb} sd = {sd} nf = {nf}
* + deltox = 0.3*(sw_tox_lv_corner - sw_tox_lv_nom) + sw_tox_lv_mc + sw_mm_tox_lv * mismatch_factor*MC_MM_SWITCH*AGAUSS(0,1.0,1)/sqrt(l*w*mult)
* + mulu0  = sw_u0_sky130_fd_pr__pfet_01v8_lvt
+ delvto = {(sw_vth0_sky130_fd_pr__pfet_01v8_lvt+sw_vth0_sky130_fd_pr__pfet_01v8_lvt_mc)*(0.005*8/l+0.995)*(0.008*7/w+0.992)*(0.0006*56/(w*l)+0.9994)+sw_mm_vth0_sky130_fd_pr__pfet_01v8_lvt*mismatch_factor*MC_MM_SWITCH*AGAUSS(0,1.0,1)/sqrt(l*w*mult)+sw_vth0_sky130_fd_pr__pfet_01v8_lvt_mc}



.model plowvt_model.1 pmos
+ level = 54 lmin = 8E-6 lmax = 2.02E-5 wmin = 7E-6
+ wmax = 1.01E-3 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 4.23E-9
+ toxm = 4.23E-9 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 9.999999999999999E22 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {7.476E-9+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {2.8E-9-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = -7.916E-9 dwb = 0 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = -0.452509 k1 = 0.64774
+ k2 = -0.04782713 k3 = 3.39 k3b = 1
+ w0 = 1E-8 lpe0 = 0 lpeb = 0
+ vbm = -3 dvtp0 = 0 dvtp1 = 0
+ dvt0 = 2.4422 dvt1 = 0.16136 dvt2 = 0.026237
+ dvt0w = 0.5 dvt1w = 1.9281E6 dvt2w = -0.032
+ vfbsdoff = 0 u0 = 2.5322839E-3 ua = -3.0054E-9
+ ub = 3.0419E-18 uc = 4.9353E-11 ud = 0
+ up = 0 lp = 1 eu = 1.67
+ vsat = 1.2376E5 a0 = 1.75209 ags = 0.385036
+ b0 = 0 b1 = 2.1073E-24 keta = -0.01258
+ a1 = 0 a2 = 0.46703705 rdsw = 484.7
+ rdswmin = 0 rdw = 0 rdwmin = 0
+ rsw = 0 rswmin = 0 prwb = 0.1
+ prwg = 0.052 wr = 1 voff = -0.1819
+ voffl = 0 minv = 0 nfactor = 2.5373
+ eta0 = 0.2 etab = -2.5E-4 dsub = 1
+ cit = -6.393105E-11 cdsc = 2.8125E-7 cdscb = 1E-4
+ cdscd = 1E-10 pclm = 0.030097 pdiblc1 = 0
+ pdiblc2 = 1.8466E-3 pdiblcb = -0.025 drout = 0.43496
+ pscbe1 = 8E8 pscbe2 = 8.6797E-9 pvag = 0
+ delta = 0.01363 fprout = 0 pdits = 0
+ pditsl = 0 pditsd = 0 lambda = 0
+ vtl = 0 lc = 5E-9 xn = 3
+ alpha0 = 5.0449517E-13 alpha1 = -4.0583656E-18 beta0 = 6.2016506
+ aigbacc = 0.43 bigbacc = 0.054 cigbacc = 0.075
+ nigbacc = 1 aigbinv = 0.35 bigbinv = 0.03
+ cigbinv = 6E-3 eigbinv = 1.1 nigbinv = 3
+ aigc = 0.43 bigc = 0.054 cigc = 0.075
+ aigsd = 0.43 bigsd = 0.054 cigsd = 0.075
+ dlcig = 0 nigc = 1 poxedge = 1
+ pigcd = 1 ntox = 1 toxref = 4.23E-9
+ agidl = 0 bgidl = 2.3E9 cgidl = 0.5
+ egidl = 0.8 noia = 3E41 noib = 0
+ noic = 0 em = 4.1E7 af = 1
+ ef = 0.88 kf = 0 lintnoi = 0
+ tnoia = 2.5E7 tnoib = 0 ntnoi = 1
+ rnoia = 0.69 rnoib = 0.34 xpart = 0
+ cgso = {2E-11/sw_func_tox_lv_ratio} cgdo = {2E-11/sw_func_tox_lv_ratio} cgbo = {1E-13/sw_func_tox_lv_ratio}
+ ckappas = 0.6 cf = 0 clc = 7E-8
+ cle = 0.492 dlc = -1.2E-8 dwc = 0
+ vfbcv = -1 noff = 2.6123 voffcv = 0.112
+ acde = 0.44 moin = 8.7 cgsl = {0/sw_func_tox_lv_ratio}
+ cgdl = {0/sw_func_tox_lv_ratio} ijthsrev = 0.1 ijthsfwd = 0.1
+ xjbvs = 1 bvs = 12.69 jss = 2.1483E-5
+ jsws = 1.4472E-10 cjs = {7.682E-04*sw_func_psd_nw_cj} mjs = 0.3362
+ mjsws = 0.2659 cjsws = {9.160236799999998E-11*sw_func_psd_nw_cj} cjswgs = {2.39155046E-10*sw_func_psd_nw_cj}
+ mjswgs = 0.9274 pbs = 0.6587 pbsws = 0.7418
+ pbswgs = 1.4338 xrcrg1 = 12 xrcrg2 = 1
+ rbpb = 50 rbpd = 50 rbps = 50
+ rbdb = 50 rbsb = 50 gbmin = 1E-12
+ tnom = 30 ute = -0.22271 kt1 = -0.60135
+ kt1l = 0 kt2 = -0.055045 ua1 = 6.8217E-10
+ ub1 = -1.4864E-19 uc1 = -9.961E-12 at = 2.856E5
+ prt = 0 njs = 1.3632 xtis = 5.2
+ tpb = 1.671E-3 tpbsw = 1.246E-3 tpbswg = 0
+ tcj = 1.2407E-3 tcjsw = 3.7357E-4 tcjswg = 2E-12
+ tvoff = 0 tvfbsdoff = 0 saref = 3E-6
+ sbref = 3E-6 wlod = 0 ku0 = 5.9E-8
+ kvsat = 0 kvth0 = 1.76E-8 tku0 = 0
+ llodku0 = 0 wlodku0 = 1 llodvth = 0
+ wlodvth = 1 lku0 = 0 wku0 = 0
+ pku0 = 0 lkvth0 = 0 wkvth0 = 7.3E-7
+ pkvth0 = 0 stk2 = 0 lodk2 = 1
+ steta0 = 0 lodeta0 = 1

.model plowvt_model.2 pmos
+ level = 54 lmin = 4E-6 lmax = 8E-6 wmin = 7E-6
+ wmax = 1.01E-3 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 4.23E-9
+ toxm = 4.23E-9 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 9.999999999999999E22 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {7.476E-9+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {2.8E-9-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = -7.916E-9 dwb = 0 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = -0.461935784 lvth0 = 7.536148200960002E-8
+ k1 = 0.64774 k2 = -0.048941198118 lk2 = 8.906306162539194E-9
+ k3 = 3.39 k3b = 1 w0 = 1E-8
+ lpe0 = 0 lpeb = 0 vbm = -3
+ dvtp0 = 0 dvtp1 = 0 dvt0 = 2.4422
+ dvt1 = 0.16136 dvt2 = 0.026237 dvt0w = 0.5
+ dvt1w = 1.9281E6 dvt2w = -0.032 vfbsdoff = 0
+ u0 = 2.45070417174E-3 lu0 = 6.521809796017425E-10 ua = -3.06421754E-9
+ lua = 4.702109417759989E-16 ub = 3.13097512E-18 lub = -7.121021393279989E-25
+ uc = 3.779220780000001E-11 luc = 9.242159716367999E-17 ud = 0
+ up = 0 lp = 1 eu = 1.67
+ vsat = 1.2376E5 a0 = 1.841424756 la0 = -7.141777733663988E-7
+ ags = 0.3685411252 lags = 1.318666271011202E-7 b0 = 0
+ b1 = 2.1073E-24 keta = -0.01258 a1 = 0
+ a2 = 0.46703705 rdsw = 484.7 rdswmin = 0
+ rdw = 0 rdwmin = 0 rsw = 0
+ rswmin = 0 prwb = 0.1 prwg = 0.052
+ wr = 1 voff = -0.1819 voffl = 0
+ minv = 0 nfactor = 2.5373 eta0 = 0.2
+ etab = -2.5E-4 dsub = 1 cit = -6.393105E-11
+ cdsc = 2.8125E-7 cdscb = 1E-4 cdscd = 1E-10
+ pclm = 0.030097 pdiblc1 = 0 pdiblc2 = 7.488388000000037E-5
+ lpdiblc2 = 1.4163807349728E-8 pdiblcb = -0.025 drout = 0.43496
+ pscbe1 = 8E8 pscbe2 = 8.6797E-9 pvag = 0
+ delta = 5.8598934E-3 ldelta = 6.211734020304E-8 fprout = 0
+ pdits = 0 pditsl = 0 pditsd = 0
+ lambda = 0 vtl = 0 lc = 5E-9
+ xn = 3 alpha0 = 5.0449517E-13 alpha1 = -4.0583656E-18
+ beta0 = 6.2016506 aigbacc = 0.43 bigbacc = 0.054
+ cigbacc = 0.075 nigbacc = 1 aigbinv = 0.35
+ bigbinv = 0.03 cigbinv = 6E-3 eigbinv = 1.1
+ nigbinv = 3 aigc = 0.43 bigc = 0.054
+ cigc = 0.075 aigsd = 0.43 bigsd = 0.054
+ cigsd = 0.075 dlcig = 0 nigc = 1
+ poxedge = 1 pigcd = 1 ntox = 1
+ toxref = 4.23E-9 agidl = 0 bgidl = 2.3E9
+ cgidl = 0.5 egidl = 0.8 noia = 3E41
+ noib = 0 noic = 0 em = 4.1E7
+ af = 1 ef = 0.88 kf = 0
+ lintnoi = 0 tnoia = 2.5E7 tnoib = 0
+ ntnoi = 1 rnoia = 0.69 rnoib = 0.34
+ xpart = 0 cgso = {2E-11/sw_func_tox_lv_ratio} cgdo = {2E-11/sw_func_tox_lv_ratio}
+ cgbo = {1E-13/sw_func_tox_lv_ratio} ckappas = 0.6 cf = 0
+ clc = 7E-8 cle = 0.492 dlc = -1.2E-8
+ dwc = 0 vfbcv = -1 noff = 2.6123
+ voffcv = 0.112 acde = 0.44 moin = 8.7
+ cgsl = {0/sw_func_tox_lv_ratio} cgdl = {0/sw_func_tox_lv_ratio} ijthsrev = 0.1
+ ijthsfwd = 0.1 xjbvs = 1 bvs = 12.69
+ jss = 2.1483E-5 jsws = 1.4472E-10 cjs = {7.682E-04*sw_func_psd_nw_cj}
+ mjs = 0.3362 mjsws = 0.2659 cjsws = {9.160236799999998E-11*sw_func_psd_nw_cj}
+ cjswgs = {2.39155046E-10*sw_func_psd_nw_cj} mjswgs = 0.9274 pbs = 0.6587
+ pbsws = 0.7418 pbswgs = 1.4338 xrcrg1 = 12
+ xrcrg2 = 1 rbpb = 50 rbpd = 50
+ rbps = 50 rbdb = 50 rbsb = 50
+ gbmin = 1E-12 tnom = 30 ute = -0.312314378
+ lute = 7.163332394831999E-7 kt1 = -0.611336 lkt1 = 7.983207840000006E-8
+ kt1l = 0 kt2 = -0.055045 ua1 = 6.68269488E-10
+ lua1 = 1.111262531327999E-16 ub1 = -1.75362536E-19 lub1 = 2.136306417984E-25
+ uc1 = -9.961E-12 at = 2.99170974E5 lat = -0.1084917945456
+ prt = 0 njs = 1.3632 xtis = 5.2
+ tpb = 1.671E-3 tpbsw = 1.246E-3 tpbswg = 0
+ tcj = 1.2407E-3 tcjsw = 3.7357E-4 tcjswg = 2E-12
+ tvoff = 0 tvfbsdoff = 0 saref = 3E-6
+ sbref = 3E-6 wlod = 0 ku0 = 5.9E-8
+ kvsat = 0 kvth0 = 1.76E-8 tku0 = 0
+ llodku0 = 0 wlodku0 = 1 llodvth = 0
+ wlodvth = 1 lku0 = 0 wku0 = 0
+ pku0 = 0 lkvth0 = 0 wkvth0 = 7.3E-7
+ pkvth0 = 0 stk2 = 0 lodk2 = 1
+ steta0 = 0 lodeta0 = 1

.model plowvt_model.3 pmos
+ level = 54 lmin = 2E-6 lmax = 4E-6 wmin = 7E-6
+ wmax = 1.01E-3 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 4.23E-9
+ toxm = 4.23E-9 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 9.999999999999999E22 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {7.476E-9+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {2.8E-9-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = -7.916E-9 dwb = 0 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = -0.4223840804 lvth0 = -8.262384285024005E-8
+ k1 = 0.64774 k2 = -0.03968662488 lk2 = -2.806016117932799E-8
+ k3 = 3.39 k3b = 1 w0 = 1E-8
+ lpe0 = 0 lpeb = 0 vbm = -3
+ dvtp0 = 0 dvtp1 = 0 dvt0 = 2.4422
+ dvt1 = 0.16136 dvt2 = 0.026237 dvt0w = 0.5
+ dvt1w = 1.9281E6 dvt2w = -0.032 vfbsdoff = 0
+ u0 = 2.32024516128E-3 lu0 = 1.173286450983169E-9 ua = -3.11313212E-9
+ lua = 6.655953401279998E-16 ub = 3.17587336E-18 lub = -8.914436691839996E-25
+ uc = 6.136577640000001E-11 luc = -1.740665252160002E-18 ud = 0
+ up = 0 lp = 1 eu = 1.67
+ vsat = 1.566795664E5 lvsat = -0.13149391602816 a0 = 2.2627309992
+ la0 = -2.397043431204481E-6 ags = 0.4230875368 lags = -8.601355939392001E-8
+ b0 = 0 b1 = 2.1073E-24 keta = -0.01258
+ a1 = 0 a2 = 0.46703705 rdsw = 484.7
+ rdswmin = 0 rdw = 0 rdwmin = 0
+ rsw = 0 rswmin = 0 prwb = 0.1
+ prwg = 0.052 wr = 1 voff = -0.1819
+ voffl = 0 minv = 0 nfactor = 2.5373
+ eta0 = 0.2 etab = -2.5E-4 dsub = 1
+ cit = -6.393105E-11 cdsc = 2.8125E-7 cdscb = 1E-4
+ cdscd = 1E-10 pclm = 0.030097 pdiblc1 = 0
+ pdiblc2 = 2.638259200000003E-4 lpdiblc2 = 1.3409097265152E-8 pdiblcb = -0.025
+ drout = 0.43496 pscbe1 = 8E8 pscbe2 = 8.6797E-9
+ pvag = 0 delta = 0.0196798608 ldelta = 6.914862420480005E-9
+ fprout = 0 pdits = 0 pditsl = 0
+ pditsd = 0 lambda = 0 vtl = 0
+ lc = 5E-9 xn = 3 alpha0 = 5.0449517E-13
+ alpha1 = -4.0583656E-18 beta0 = 6.2016506 aigbacc = 0.43
+ bigbacc = 0.054 cigbacc = 0.075 nigbacc = 1
+ aigbinv = 0.35 bigbinv = 0.03 cigbinv = 6E-3
+ eigbinv = 1.1 nigbinv = 3 aigc = 0.43
+ bigc = 0.054 cigc = 0.075 aigsd = 0.43
+ bigsd = 0.054 cigsd = 0.075 dlcig = 0
+ nigc = 1 poxedge = 1 pigcd = 1
+ ntox = 1 toxref = 4.23E-9 agidl = 0
+ bgidl = 2.3E9 cgidl = 0.5 egidl = 0.8
+ noia = 3E41 noib = 0 noic = 0
+ em = 4.1E7 af = 1 ef = 0.88
+ kf = 0 lintnoi = 0 tnoia = 2.5E7
+ tnoib = 0 ntnoi = 1 rnoia = 0.69
+ rnoib = 0.34 xpart = 0 cgso = {2E-11/sw_func_tox_lv_ratio}
+ cgdo = {2E-11/sw_func_tox_lv_ratio} cgbo = {1E-13/sw_func_tox_lv_ratio} ckappas = 0.6
+ cf = 0 clc = 7E-8 cle = 0.492
+ dlc = -1.2E-8 dwc = 0 vfbcv = -1
+ noff = 2.6123 voffcv = 0.112 acde = 0.44
+ moin = 8.7 cgsl = {0/sw_func_tox_lv_ratio} cgdl = {0/sw_func_tox_lv_ratio}
+ ijthsrev = 0.1 ijthsfwd = 0.1 xjbvs = 1
+ bvs = 12.69 jss = 2.1483E-5 jsws = 1.4472E-10
+ cjs = {7.682E-04*sw_func_psd_nw_cj} mjs = 0.3362 mjsws = 0.2659
+ cjsws = {9.160236799999998E-11*sw_func_psd_nw_cj} cjswgs = {2.39155046E-10*sw_func_psd_nw_cj} mjswgs = 0.9274
+ pbs = 0.6587 pbsws = 0.7418 pbswgs = 1.4338
+ xrcrg1 = 12 xrcrg2 = 1 rbpb = 50
+ rbpd = 50 rbps = 50 rbdb = 50
+ rbsb = 50 gbmin = 1E-12 tnom = 30
+ ute = -0.13298 kt1 = -0.59135 kt1l = 0
+ kt2 = -0.055045 ua1 = 6.9609E-10 ub1 = -1.57126034E-19
+ lub1 = 1.407867582096E-25 uc1 = -9.961E-12 at = 3.78032304E5
+ lat = -0.4234954910976 prt = 0 njs = 1.3632
+ xtis = 5.2 tpb = 1.671E-3 tpbsw = 1.246E-3
+ tpbswg = 0 tcj = 1.2407E-3 tcjsw = 3.7357E-4
+ tcjswg = 2E-12 tvoff = 0 tvfbsdoff = 0
+ saref = 3E-6 sbref = 3E-6 wlod = 0
+ ku0 = 5.9E-8 kvsat = 0 kvth0 = 1.76E-8
+ tku0 = 0 llodku0 = 0 wlodku0 = 1
+ llodvth = 0 wlodvth = 1 lku0 = 0
+ wku0 = 0 pku0 = 0 lkvth0 = 0
+ wkvth0 = 7.3E-7 pkvth0 = 0 stk2 = 0
+ lodk2 = 1 steta0 = 0 lodeta0 = 1

.model plowvt_model.4 pmos
+ level = 54 lmin = 1.5E-6 lmax = 2E-6 wmin = 7E-6
+ wmax = 1.01E-3 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 4.23E-9
+ toxm = 4.23E-9 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 9.999999999999999E22 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {7.476E-9+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {2.8E-9-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = -7.916E-9 dwb = 0 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = -0.4703903488 lvth0 = 1.311985884672005E-8
+ k1 = 0.64774 k2 = -0.04752564752 lk2 = -1.242601442611199E-8
+ k3 = 3.39 k3b = 1 w0 = 1E-8
+ lpe0 = 0 lpeb = 0 vbm = -3
+ dvtp0 = 0 dvtp1 = 0 dvt0 = 2.4422
+ dvt1 = 0.16136 dvt2 = 0.026237 dvt0w = 0.5
+ dvt1w = 1.9281E6 dvt2w = -0.032 vfbsdoff = 0
+ u0 = 3.15488624448E-3 lu0 = -4.913217253509119E-10 ua = -2.23484064E-9
+ lua = -1.086069187584E-15 ub = 1.831961120000001E-18 lub = 1.788854902271998E-24
+ uc = 2.748768160000001E-11 luc = 6.582580701695997E-17 ud = 0
+ up = 0 lp = 1 eu = 1.67
+ vsat = 9.0748E4 a0 = 1.1005741184 la0 = -7.923774813696E-8
+ ags = 0.167247104 lags = 4.242345997823998E-7 b0 = 0
+ b1 = 2.1073E-24 keta = -0.01258 a1 = 0
+ a2 = 0.46703705 rdsw = 484.7 rdswmin = 0
+ rdw = 0 rdwmin = 0 rsw = 0
+ rswmin = 0 prwb = 0.1 prwg = 0.052
+ wr = 1 voff = -0.1819 voffl = 0
+ minv = 0 nfactor = 2.5373 eta0 = 0.2
+ etab = -2.5E-4 dsub = 1 cit = -6.393105E-11
+ cdsc = 2.8125E-7 cdscb = 1E-4 cdscd = 1E-10
+ pclm = 0.030097 pdiblc1 = 0 pdiblc2 = -3.278730240000004E-3
+ lpdiblc2 = 2.0474371270656E-8 pdiblcb = -0.025 drout = 0.43496
+ pscbe1 = 8E8 pscbe2 = 8.6797E-9 pvag = 0
+ delta = 0.0169691504 ldelta = 1.232110324224E-8 fprout = 0
+ pdits = 0 pditsl = 0 pditsd = 0
+ lambda = 0 vtl = 0 lc = 5E-9
+ xn = 3 alpha0 = 5.0449517E-13 alpha1 = -4.0583656E-18
+ beta0 = 6.2016506 aigbacc = 0.43 bigbacc = 0.054
+ cigbacc = 0.075 nigbacc = 1 aigbinv = 0.35
+ bigbinv = 0.03 cigbinv = 6E-3 eigbinv = 1.1
+ nigbinv = 3 aigc = 0.43 bigc = 0.054
+ cigc = 0.075 aigsd = 0.43 bigsd = 0.054
+ cigsd = 0.075 dlcig = 0 nigc = 1
+ poxedge = 1 pigcd = 1 ntox = 1
+ toxref = 4.23E-9 agidl = 0 bgidl = 2.3E9
+ cgidl = 0.5 egidl = 0.8 noia = 3E41
+ noib = 0 noic = 0 em = 4.1E7
+ af = 1 ef = 0.88 kf = 0
+ lintnoi = 0 tnoia = 2.5E7 tnoib = 0
+ ntnoi = 1 rnoia = 0.69 rnoib = 0.34
+ xpart = 0 cgso = {2E-11/sw_func_tox_lv_ratio} cgdo = {2E-11/sw_func_tox_lv_ratio}
+ cgbo = {1E-13/sw_func_tox_lv_ratio} ckappas = 0.6 cf = 0
+ clc = 7E-8 cle = 0.492 dlc = -1.2E-8
+ dwc = 0 vfbcv = -1 noff = 2.6123
+ voffcv = 0.112 acde = 0.44 moin = 8.7
+ cgsl = {0/sw_func_tox_lv_ratio} cgdl = {0/sw_func_tox_lv_ratio} ijthsrev = 0.1
+ ijthsfwd = 0.1 xjbvs = 1 bvs = 12.69
+ jss = 2.1483E-5 jsws = 1.4472E-10 cjs = {7.682E-04*sw_func_psd_nw_cj}
+ mjs = 0.3362 mjsws = 0.2659 cjsws = {9.160236799999998E-11*sw_func_psd_nw_cj}
+ cjswgs = {2.39155046E-10*sw_func_psd_nw_cj} mjswgs = 0.9274 pbs = 0.6587
+ pbsws = 0.7418 pbswgs = 1.4338 xrcrg1 = 12
+ xrcrg2 = 1 rbpb = 50 rbpd = 50
+ rbps = 50 rbdb = 50 rbsb = 50
+ gbmin = 1E-12 tnom = 30 ute = -0.13298
+ kt1 = -0.59135 kt1l = 0 kt2 = -0.055045
+ ua1 = 8.001002400000001E-10 lua1 = -2.074380226560002E-16 ub1 = -3.12473336E-19
+ lub1 = 4.506114173184001E-25 uc1 = -9.961E-12 at = 2.05829584E5
+ lat = -0.0800543863296 prt = 0 njs = 1.3632
+ xtis = 5.2 tpb = 1.671E-3 tpbsw = 1.246E-3
+ tpbswg = 0 tcj = 1.2407E-3 tcjsw = 3.7357E-4
+ tcjswg = 2E-12 tvoff = 0 tvfbsdoff = 0
+ saref = 3E-6 sbref = 3E-6 wlod = 0
+ ku0 = 5.9E-8 kvsat = 0 kvth0 = 1.76E-8
+ tku0 = 0 llodku0 = 0 wlodku0 = 1
+ llodvth = 0 wlodvth = 1 lku0 = 0
+ wku0 = 0 pku0 = 0 lkvth0 = 0
+ wkvth0 = 7.3E-7 pkvth0 = 0 stk2 = 0
+ lodk2 = 1 steta0 = 0 lodeta0 = 1

.model plowvt_model.5 pmos
+ level = 54 lmin = 1E-6 lmax = 1.5E-6 wmin = 7E-6
+ wmax = 1.01E-3 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 4.23E-9
+ toxm = 4.23E-9 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 9.999999999999999E22 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {7.476E-9+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {2.8E-9-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = -7.916E-9 dwb = 0 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = -0.4490338288 lvth0 = -1.879532464127999E-8
+ k1 = 0.64774 k2 = -0.05110258288 lk2 = -7.080642224128E-9
+ k3 = 3.39 k3b = 1 w0 = 1E-8
+ lpe0 = 0 lpeb = 0 vbm = -3
+ dvtp0 = 0 dvtp1 = 0 dvt0 = 2.4422
+ dvt1 = 0.16136 dvt2 = 0.026237 dvt0w = 0.5
+ dvt1w = 1.9281E6 dvt2w = -0.032 vfbsdoff = 0
+ u0 = 2.0291928736E-3 lu0 = 1.19091444809216E-9 ua = -3.153121440000001E-9
+ lua = 2.862096399360005E-16 ub = 3.14096944E-18 lub = -1.673271311359996E-25
+ uc = 6.93721856E-11 luc = 3.233604239360006E-18 ud = 0
+ up = 0 lp = 1 eu = 1.67
+ vsat = 9.00260656E4 lvsat = 1.07885876736E-3 a0 = 0.8695573776
+ la0 = 2.659936693145603E-7 ags = -0.021289552 lags = 7.059837785088002E-7
+ b0 = 0 b1 = 2.1073E-24 keta = -0.01258
+ a1 = 0 a2 = 0.46703705 rdsw = 484.7
+ rdswmin = 0 rdw = 0 rdwmin = 0
+ rsw = 0 rswmin = 0 prwb = 0.1
+ prwg = 0.052 wr = 1 voff = -0.15296296
+ lvoff = -4.324351257600003E-8 voffl = 0 minv = 0
+ nfactor = 2.59775952 lnfactor = -9.035070668800062E-8 eta0 = 0.2
+ etab = -2.5E-4 dsub = 1 cit = -6.393105E-11
+ cdsc = 2.8125E-7 cdscb = 1E-4 cdscd = 1E-10
+ pclm = 0.030097 pdiblc1 = 0 pdiblc2 = 5.973279999999994E-4
+ lpdiblc2 = 1.46819898368E-8 pdiblcb = -0.025 drout = 0.43496
+ pscbe1 = 8E8 pscbe2 = 8.6797E-9 pvag = 0
+ delta = 0.0102363472 ldelta = 2.238260434432001E-8 fprout = 0
+ pdits = 0 pditsl = 0 pditsd = 0
+ lambda = 0 vtl = 0 lc = 5E-9
+ xn = 3 alpha0 = 5.0449517E-13 alpha1 = -4.0583656E-18
+ beta0 = 6.2016506 aigbacc = 0.43 bigbacc = 0.054
+ cigbacc = 0.075 nigbacc = 1 aigbinv = 0.35
+ bigbinv = 0.03 cigbinv = 6E-3 eigbinv = 1.1
+ nigbinv = 3 aigc = 0.43 bigc = 0.054
+ cigc = 0.075 aigsd = 0.43 bigsd = 0.054
+ cigsd = 0.075 dlcig = 0 nigc = 1
+ poxedge = 1 pigcd = 1 ntox = 1
+ toxref = 4.23E-9 agidl = 0 bgidl = 2.3E9
+ cgidl = 0.5 egidl = 0.8 noia = 3E41
+ noib = 0 noic = 0 em = 4.1E7
+ af = 1 ef = 0.88 kf = 0
+ lintnoi = 0 tnoia = 2.5E7 tnoib = 0
+ ntnoi = 1 rnoia = 0.69 rnoib = 0.34
+ xpart = 0 cgso = {2E-11/sw_func_tox_lv_ratio} cgdo = {2E-11/sw_func_tox_lv_ratio}
+ cgbo = {1E-13/sw_func_tox_lv_ratio} ckappas = 0.6 cf = 0
+ clc = 7E-8 cle = 0.492 dlc = -1.2E-8
+ dwc = 0 vfbcv = -1 noff = 2.6123
+ voffcv = 0.112 acde = 0.44 moin = 8.7
+ cgsl = {0/sw_func_tox_lv_ratio} cgdl = {0/sw_func_tox_lv_ratio} ijthsrev = 0.1
+ ijthsfwd = 0.1 xjbvs = 1 bvs = 12.69
+ jss = 2.1483E-5 jsws = 1.4472E-10 cjs = {7.682E-04*sw_func_psd_nw_cj}
+ mjs = 0.3362 mjsws = 0.2659 cjsws = {9.160236799999998E-11*sw_func_psd_nw_cj}
+ cjswgs = {2.39155046E-10*sw_func_psd_nw_cj} mjswgs = 0.9274 pbs = 0.6587
+ pbsws = 0.7418 pbswgs = 1.4338 xrcrg1 = 12
+ xrcrg2 = 1 rbpb = 50 rbpd = 50
+ rbps = 50 rbdb = 50 rbsb = 50
+ gbmin = 1E-12 tnom = 30 ute = 0.05615488
+ lute = -2.826431646720001E-7 kt1 = -0.651014 lkt1 = 8.91618816000001E-8
+ kt1l = 0 kt2 = -0.0933612208 lkt2 = 5.725976036352E-8
+ ua1 = 6.6129E-10 ub1 = -1.05044528E-20 lub1 = -6.508817356799988E-28
+ uc1 = -9.961E-12 at = 2.04346672E5 lat = -0.0778383226368
+ prt = 0 njs = 1.3632 xtis = 5.2
+ tpb = 1.671E-3 tpbsw = 1.246E-3 tpbswg = 0
+ tcj = 1.2407E-3 tcjsw = 3.7357E-4 tcjswg = 2E-12
+ tvoff = 0 tvfbsdoff = 0 saref = 3E-6
+ sbref = 3E-6 wlod = 0 ku0 = 5.9E-8
+ kvsat = 0 kvth0 = 1.76E-8 tku0 = 0
+ llodku0 = 0 wlodku0 = 1 llodvth = 0
+ wlodvth = 1 lku0 = 0 wku0 = 0
+ pku0 = 0 lkvth0 = 0 wkvth0 = 7.3E-7
+ pkvth0 = 0 stk2 = 0 lodk2 = 1
+ steta0 = 0 lodeta0 = 1

.model plowvt_model.6 pmos
+ level = 54 lmin = 5E-7 lmax = 1E-6 wmin = 7E-6
+ wmax = 1.01E-3 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 4.23E-9
+ toxm = 4.23E-9 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 9.999999999999999E22 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {7.476E-9+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {2.8E-9-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = -7.916E-9 dwb = 0 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = -0.4731173008 lvth0 = 5.153279915519995E-9
+ k1 = 0.64774 k2 = -0.06360790704 lk2 = 5.354652120576E-9
+ k3 = 3.39 k3b = 1 w0 = 1E-8
+ lpe0 = 0 lpeb = 0 vbm = -3
+ dvtp0 = 0 dvtp1 = 0 dvt0 = 2.4422
+ dvt1 = 0.16136 dvt2 = 0.026237 dvt0w = 0.5
+ dvt1w = 1.9281E6 dvt2w = -0.032 vfbsdoff = 0
+ u0 = 3.2439924224E-3 lu0 = -1.708222323456021E-11 ua = -2.78985456E-9
+ lua = -7.502294553599983E-17 ub = 2.82507216E-18 lub = 1.46801124096E-25
+ uc = 7.576047360000001E-11 luc = -3.118909347840004E-18 ud = 0
+ up = 0 lp = 1 eu = 1.67
+ vsat = 6.32733136E4 lvsat = 0.02768179535616 a0 = 1.2056064592
+ la0 = -6.817353742848001E-8 ags = 0.95347064 lags = -2.63317756416E-7
+ b0 = 7.305551039999999E-7 lb0 = -7.264639954176E-13 b1 = 2.1073E-24
+ keta = -0.01258 a1 = 0 a2 = 0.46703705
+ rdsw = 484.7 rdswmin = 0 rdw = 0
+ rdwmin = 0 rsw = 0 rswmin = 0
+ prwb = 0.1 prwg = 0.052 wr = 1
+ voff = -0.21083704 lvoff = 1.430647257600001E-8 voffl = 0
+ minv = 0 nfactor = 2.47684048 lnfactor = 2.98911866880002E-8
+ eta0 = 0.2 etab = -2.5E-4 dsub = 1
+ cit = -6.393105E-11 cdsc = 2.8125E-7 cdscb = 1E-4
+ cdscd = 1E-10 pclm = 0.030097 pdiblc1 = 0
+ pdiblc2 = -0.0227473408 lpdiblc2 = 3.789592849152E-8 pdiblcb = -0.025
+ drout = 0.43496 pscbe1 = 8E8 pscbe2 = 8.6797E-9
+ pvag = 0 delta = 0.021368856 ldelta = 1.131243759359999E-8
+ fprout = 0 pdits = 0 pditsl = 0
+ pditsd = 0 lambda = 0 vtl = 0
+ lc = 5E-9 xn = 3 alpha0 = 5.0449517E-13
+ alpha1 = -4.0583656E-18 beta0 = 6.2016506 aigbacc = 0.43
+ bigbacc = 0.054 cigbacc = 0.075 nigbacc = 1
+ aigbinv = 0.35 bigbinv = 0.03 cigbinv = 6E-3
+ eigbinv = 1.1 nigbinv = 3 aigc = 0.43
+ bigc = 0.054 cigc = 0.075 aigsd = 0.43
+ bigsd = 0.054 cigsd = 0.075 dlcig = 0
+ nigc = 1 poxedge = 1 pigcd = 1
+ ntox = 1 toxref = 4.23E-9 agidl = 0
+ bgidl = 2.3E9 cgidl = 0.5 egidl = 0.8
+ noia = 3E41 noib = 0 noic = 0
+ em = 4.1E7 af = 1 ef = 0.88
+ kf = 0 lintnoi = 0 tnoia = 2.5E7
+ tnoib = 0 ntnoi = 1 rnoia = 0.69
+ rnoib = 0.34 xpart = 0 cgso = {2E-11/sw_func_tox_lv_ratio}
+ cgdo = {2E-11/sw_func_tox_lv_ratio} cgbo = {1E-13/sw_func_tox_lv_ratio} ckappas = 0.6
+ cf = 0 clc = 7E-8 cle = 0.492
+ dlc = -1.2E-8 dwc = 0 vfbcv = -1
+ noff = 2.6123 voffcv = 0.112 acde = 0.44
+ moin = 8.7 cgsl = {0/sw_func_tox_lv_ratio} cgdl = {0/sw_func_tox_lv_ratio}
+ ijthsrev = 0.1 ijthsfwd = 0.1 xjbvs = 1
+ bvs = 12.69 jss = 2.1483E-5 jsws = 1.4472E-10
+ cjs = {7.682E-04*sw_func_psd_nw_cj} mjs = 0.3362 mjsws = 0.2659
+ cjsws = {9.160236799999998E-11*sw_func_psd_nw_cj} cjswgs = {2.39155046E-10*sw_func_psd_nw_cj} mjswgs = 0.9274
+ pbs = 0.6587 pbsws = 0.7418 pbswgs = 1.4338
+ xrcrg1 = 12 xrcrg2 = 1 rbpb = 50
+ rbpd = 50 rbps = 50 rbdb = 50
+ rbsb = 50 gbmin = 1E-12 tnom = 30
+ ute = -0.05958848 lute = -1.67547967488E-7 kt1 = -0.491530832
+ lkt1 = -6.942818065919995E-8 kt1l = 0 kt2 = -0.0157696432
+ lkt2 = -1.989730440192E-8 ua1 = 4.28862672E-10 lua1 = 2.311257349632E-16
+ ub1 = 5.703157168E-19 lub1 = -5.7821845838592E-25 uc1 = -2.284941472E-11
+ luc1 = 1.2816239597568E-17 at = 1.920565792E5 lat = -0.06561705435648
+ prt = 0 njs = 1.3632 xtis = 5.2
+ tpb = 1.671E-3 tpbsw = 1.246E-3 tpbswg = 0
+ tcj = 1.2407E-3 tcjsw = 3.7357E-4 tcjswg = 2E-12
+ tvoff = 0 tvfbsdoff = 0 saref = 2.74E-6
+ sbref = 2.74E-6 wlod = 0 ku0 = 5.9E-8
+ kvsat = 0 kvth0 = 1.76E-8 tku0 = 0
+ llodku0 = 0 wlodku0 = 1 llodvth = 0
+ wlodvth = 1 lku0 = 0 wku0 = 0
+ pku0 = 0 lkvth0 = 0 wkvth0 = 7.3E-7
+ pkvth0 = 0 stk2 = 0 lodk2 = 1
+ steta0 = 0 lodeta0 = 1

.model plowvt_model.7 pmos
+ level = 54 lmin = 3.5E-7 lmax = 5E-7 wmin = 7E-6
+ wmax = 1.01E-3 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 4.23E-9
+ toxm = 4.23E-9 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 9.999999999999999E22 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {7.476E-9+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {2.8E-9-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = -7.916E-9 dwb = 0 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = -0.479241272 lvth0 = 8.180971276800022E-9
+ k1 = 0.64774 k2 = -0.0662396664 lk2 = 6.655793948159998E-9
+ k3 = 3.39 k3b = 1 w0 = 1E-8
+ lpe0 = 0 lpeb = 0 vbm = -3
+ dvtp0 = 0 dvtp1 = 0 dvt0 = 2.4422
+ dvt1 = 0.16136 dvt2 = 0.026237 dvt0w = 0.5
+ dvt1w = 1.9281E6 dvt2w = -0.032 vfbsdoff = 0
+ u0 = 2.40470448E-3 lu0 = 3.978617354880002E-10 ua = -3.0740792E-9
+ lua = 6.54977164799999E-17 ub = 3.03016E-18 lub = 4.540569599999976E-26
+ uc = 8.394894399999999E-11 luc = -7.167289113599997E-18 ud = 0
+ up = 0 lp = 1 eu = 1.67
+ vsat = 1.58275336E5 lvsat = -0.0192872045184 a0 = 1.22318864
+ la0 = -7.686616761599996E-8 ags = 0.411112 lags = 4.824355199999972E-9
+ b0 = -2.43518368E-6 lb0 = 8.38677259392E-13 b1 = 2.1073E-24
+ keta = -0.01258 a1 = 0 a2 = 0.46703705
+ rdsw = 484.7 rdswmin = 0 rdw = 0
+ rdwmin = 0 rsw = 0 rswmin = 0
+ prwb = 0.1 prwg = 0.052 wr = 1
+ voff = -0.1819 voffl = 0 minv = 0
+ nfactor = 2.5373 eta0 = 0.2 etab = -2.5E-4
+ dsub = 1 cit = -6.393105E-11 cdsc = 2.8125E-7
+ cdscb = 1E-4 cdscd = 1E-10 pclm = 0.030097
+ pdiblc1 = 0 pdiblc2 = -0.088488032 lpdiblc2 = 7.03981262208E-8
+ pdiblcb = -0.025 drout = 0.43496 pscbe1 = 8E8
+ pscbe2 = 8.6797E-9 pvag = 0 delta = 0.024897016
+ ldelta = 9.5681152896E-9 fprout = 0 pdits = 0
+ pditsl = 0 pditsd = 0 lambda = 0
+ vtl = 0 lc = 5E-9 xn = 3
+ alpha0 = 5.0449517E-13 alpha1 = -4.0583656E-18 beta0 = 6.2016506
+ aigbacc = 0.43 bigbacc = 0.054 cigbacc = 0.075
+ nigbacc = 1 aigbinv = 0.35 bigbinv = 0.03
+ cigbinv = 6E-3 eigbinv = 1.1 nigbinv = 3
+ aigc = 0.43 bigc = 0.054 cigc = 0.075
+ aigsd = 0.43 bigsd = 0.054 cigsd = 0.075
+ dlcig = 0 nigc = 1 poxedge = 1
+ pigcd = 1 ntox = 1 toxref = 4.23E-9
+ agidl = 0 bgidl = 2.3E9 cgidl = 0.5
+ egidl = 0.8 noia = 3E41 noib = 0
+ noic = 0 em = 4.1E7 af = 1
+ ef = 0.88 kf = 0 lintnoi = 0
+ tnoia = 2.5E7 tnoib = 0 ntnoi = 1
+ rnoia = 0.69 rnoib = 0.34 xpart = 0
+ cgso = {2E-11/sw_func_tox_lv_ratio} cgdo = {2E-11/sw_func_tox_lv_ratio} cgbo = {1E-13/sw_func_tox_lv_ratio}
+ ckappas = 0.6 cf = 0 clc = 7E-8
+ cle = 0.492 dlc = -1.2E-8 dwc = 0
+ vfbcv = -1 noff = 2.6123 voffcv = 0.112
+ acde = 0.44 moin = 8.7 cgsl = {0/sw_func_tox_lv_ratio}
+ cgdl = {0/sw_func_tox_lv_ratio} ijthsrev = 0.1 ijthsfwd = 0.1
+ xjbvs = 1 bvs = 12.69 jss = 2.1483E-5
+ jsws = 1.4472E-10 cjs = {7.682E-04*sw_func_psd_nw_cj} mjs = 0.3362
+ mjsws = 0.2659 cjsws = {9.160236799999998E-11*sw_func_psd_nw_cj} cjswgs = {2.39155046E-10*sw_func_psd_nw_cj}
+ mjswgs = 0.9274 pbs = 0.6587 pbsws = 0.7418
+ pbswgs = 1.4338 xrcrg1 = 12 xrcrg2 = 1
+ rbpb = 50 rbpd = 50 rbps = 50
+ rbdb = 50 rbsb = 50 gbmin = 1E-12
+ tnom = 30 ute = -0.39848 kt1 = -0.65492
+ lkt1 = 1.135142400000001E-8 kt1l = 0 kt2 = -0.056015
+ ua1 = 8.9635E-10 ub1 = -5.9922E-19 uc1 = 3.0734E-12
+ at = 1.37677816E5 lat = -0.0387321938304 prt = 0
+ njs = 1.3632 xtis = 5.2 tpb = 1.671E-3
+ tpbsw = 1.246E-3 tpbswg = 0 tcj = 1.2407E-3
+ tcjsw = 3.7357E-4 tcjswg = 2E-12 tvoff = 0
+ tvfbsdoff = 0 saref = 1.74E-6 sbref = 1.74E-6
+ wlod = 0 ku0 = 5.9E-8 kvsat = 0
+ kvth0 = 1.76E-8 tku0 = 0 llodku0 = 0
+ wlodku0 = 1 llodvth = 0 wlodvth = 1
+ lku0 = 0 wku0 = 0 pku0 = 0
+ lkvth0 = 0 wkvth0 = 7.3E-7 pkvth0 = 0
+ stk2 = 0 lodk2 = 1 steta0 = 0
+ lodeta0 = 1

.model plowvt_model.8 pmos
+ level = 54 lmin = 8E-6 lmax = 2.02E-5 wmin = 5E-6
+ wmax = 7E-6 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 4.23E-9
+ toxm = 4.23E-9 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 9.999999999999999E22 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {7.476E-9+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {2.8E-9-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = -7.916E-9 dwb = 0 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = -0.486529460076 wvth0 = 2.37634546612944E-7
+ k1 = 0.64774 k2 = -0.05280901249452 wk2 = 3.479868835458201E-8
+ k3 = 3.39 k3b = 1 w0 = 1E-8
+ lpe0 = 0 lpeb = 0 vbm = -3
+ dvtp0 = 0 dvtp1 = 0 dvt0 = 2.4422
+ dvt1 = 0.16136 dvt2 = 0.026237 dvt0w = 0.5
+ dvt1w = 1.9281E6 dvt2w = -0.032 vfbsdoff = 0
+ u0 = 2.6027896771356E-3 wu0 = -4.924862375694697E-10 ua = -3.1218008708E-9
+ wua = 8.130656697797957E-16 ub = 3.2320795812E-18 wub = -1.3284135033019E-24
+ uc = 5.087094711600001E-11 wuc = -1.060293346672162E-17 ud = 0
+ up = 0 lp = 1 eu = 1.67
+ vsat = 1.2376E5 a0 = 1.74665629768 wa0 = 3.795467152291259E-8
+ ags = 0.437022573068 wags = -3.631287082354875E-7 b0 = 0
+ b1 = 2.1073E-24 keta = -0.01258 a1 = 0
+ a2 = 0.46703705 rdsw = 484.7 rdswmin = 0
+ rdw = 0 rdwmin = 0 rsw = 0
+ rswmin = 0 prwb = 0.1 prwg = 0.052
+ wr = 1 voff = -0.1819 voffl = 0
+ minv = 0 nfactor = 2.5373 eta0 = 0.2
+ etab = -2.5E-4 dsub = 1 cit = -6.393105E-11
+ cdsc = 2.8125E-7 cdscb = 1E-4 cdscd = 1E-10
+ pclm = 0.030097 pdiblc1 = 0 pdiblc2 = 2.3508376052E-3
+ wpdiblc2 = -3.522123875727051E-9 pdiblcb = -0.025 drout = 0.43496
+ pscbe1 = 8E8 pscbe2 = 8.6797E-9 pvag = 0
+ delta = 3.48542732E-3 wdelta = 7.086032710928865E-8 fprout = 0
+ pdits = 0 pditsl = 0 pditsd = 0
+ lambda = 0 vtl = 0 lc = 5E-9
+ xn = 3 alpha0 = 5.0449517E-13 alpha1 = -4.0583656E-18
+ beta0 = 6.2016506 aigbacc = 0.43 bigbacc = 0.054
+ cigbacc = 0.075 nigbacc = 1 aigbinv = 0.35
+ bigbinv = 0.03 cigbinv = 6E-3 eigbinv = 1.1
+ nigbinv = 3 aigc = 0.43 bigc = 0.054
+ cigc = 0.075 aigsd = 0.43 bigsd = 0.054
+ cigsd = 0.075 dlcig = 0 nigc = 1
+ poxedge = 1 pigcd = 1 ntox = 1
+ toxref = 4.23E-9 agidl = 0 bgidl = 2.3E9
+ cgidl = 0.5 egidl = 0.8 noia = 3E41
+ noib = 0 noic = 0 em = 4.1E7
+ af = 1 ef = 0.88 kf = 0
+ lintnoi = 0 tnoia = 2.5E7 tnoib = 0
+ ntnoi = 1 rnoia = 0.69 rnoib = 0.34
+ xpart = 0 cgso = {2E-11/sw_func_tox_lv_ratio} cgdo = {2E-11/sw_func_tox_lv_ratio}
+ cgbo = {1E-13/sw_func_tox_lv_ratio} ckappas = 0.6 cf = 0
+ clc = 7E-8 cle = 0.492 dlc = -1.2E-8
+ dwc = 0 vfbcv = -1 noff = 2.6123
+ voffcv = 0.112 acde = 0.44 moin = 8.7
+ cgsl = {0/sw_func_tox_lv_ratio} cgdl = {0/sw_func_tox_lv_ratio} ijthsrev = 0.1
+ ijthsfwd = 0.1 xjbvs = 1 bvs = 12.69
+ jss = 2.1483E-5 jsws = 1.4472E-10 cjs = {7.682E-04*sw_func_psd_nw_cj}
+ mjs = 0.3362 mjsws = 0.2659 cjsws = {9.160236799999998E-11*sw_func_psd_nw_cj}
+ cjswgs = {2.39155046E-10*sw_func_psd_nw_cj} mjswgs = 0.9274 pbs = 0.6587
+ pbsws = 0.7418 pbswgs = 1.4338 xrcrg1 = 12
+ xrcrg2 = 1 rbpb = 50 rbpd = 50
+ rbps = 50 rbdb = 50 rbsb = 50
+ gbmin = 1E-12 tnom = 30 ute = -0.22271
+ kt1 = -0.60135 kt1l = 0 kt2 = -0.055045
+ ua1 = 6.8217E-10 ub1 = -1.4864E-19 uc1 = -9.961E-12
+ at = 2.856E5 prt = 0 njs = 1.3632
+ xtis = 5.2 tpb = 1.671E-3 tpbsw = 1.246E-3
+ tpbswg = 0 tcj = 1.2407E-3 tcjsw = 3.7357E-4
+ tcjswg = 2E-12 tvoff = 0 tvfbsdoff = 0
+ saref = 3E-6 sbref = 3E-6 wlod = 0
+ ku0 = 5.9E-8 kvsat = 0 kvth0 = 1.76E-8
+ tku0 = 0 llodku0 = 0 wlodku0 = 1
+ llodvth = 0 wlodvth = 1 lku0 = 0
+ wku0 = 0 pku0 = 0 lkvth0 = 0
+ wkvth0 = 7.3E-7 pkvth0 = 0 stk2 = 0
+ lodk2 = 1 steta0 = 0 lodeta0 = 1

.model plowvt_model.9 pmos
+ level = 54 lmin = 4E-6 lmax = 8E-6 wmin = 5E-6
+ wmax = 7E-6 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 4.23E-9
+ toxm = 4.23E-9 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 9.999999999999999E22 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {7.476E-9+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {2.8E-9-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = -7.916E-9 dwb = 0 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = -0.498131660199634 lvth0 = 9.27526286683773E-8
+ wvth0 = 2.528299326564993E-7 pvth0 = -1.214779941865989E-13 k1 = 0.64774
+ k2 = -0.058057192628798 lk2 = 4.195605126547001E-8 wk2 = 6.367565922565886E-8
+ pk2 = -2.308540559317367E-13 k3 = 3.39 k3b = 1
+ w0 = 1E-8 lpe0 = 0 lpeb = 0
+ vbm = -3 dvtp0 = 0 dvtp1 = 0
+ dvt0 = 2.4422 dvt1 = 0.16136 dvt2 = 0.026237
+ dvt0w = 0.5 dvt1w = 1.9281E6 dvt2w = -0.032
+ vfbsdoff = 0 u0 = 2.370302029308788E-3 lu0 = 1.858599251786666E-9
+ wu0 = 5.616128241848532E-10 pu0 = -8.426889539288758E-15 ua = -3.327222540870959E-9
+ lua = 1.642222999215279E-15 wua = 1.837102555323692E-15 pua = -8.186560477792127E-21
+ ub = 3.54317657560288E-18 lub = -2.48703381205438E-24 wub = -2.879246953055986E-24
+ pub = 1.239798293071406E-29 uc = 1.049460289848722E-11 luc = 3.227846462124842E-16
+ wuc = 1.906750805221021E-16 puc = -1.609096955032252E-21 ud = 0
+ up = 0 lp = 1 eu = 1.67
+ vsat = 1.2376E5 a0 = 2.069238473526343 la0 = -2.57885094658601E-6
+ wa0 = -1.591289751979952E-6 pa0 = 1.30248316192513E-11 ags = 0.489045839059059
+ lags = -4.158947976389233E-7 wags = -8.417312105317939E-7 pags = 3.826139844357592E-12
+ b0 = 0 b1 = 2.1073E-24 keta = -0.01258
+ a1 = 0 a2 = 0.46703705 rdsw = 484.7
+ rdswmin = 0 rdw = 0 rdwmin = 0
+ rsw = 0 rswmin = 0 prwb = 0.1
+ prwg = 0.052 wr = 1 voff = -0.1819
+ voffl = 0 minv = 0 nfactor = 2.5373
+ eta0 = 0.2 etab = -2.5E-4 dsub = 1
+ cit = -6.393105E-11 cdsc = 2.8125E-7 cdscb = 1E-4
+ cdscd = 1E-10 pclm = 0.030097 pdiblc1 = 0
+ pdiblc2 = -1.270175929176788E-4 lpdiblc2 = 1.980896559583197E-8 wpdiblc2 = 1.41029147960069E-9
+ ppdiblc2 = -3.943170131663209E-14 pdiblcb = -0.025 drout = 0.43496
+ pscbe1 = 8E8 pscbe2 = 8.6797E-9 pvag = 0
+ delta = -0.011930993160781 ldelta = 1.23245031891554E-7 wdelta = 1.242701965896088E-7
+ pdelta = -4.269798605734718E-13 fprout = 0 pdits = 0
+ pditsl = 0 pditsd = 0 lambda = 0
+ vtl = 0 lc = 5E-9 xn = 3
+ alpha0 = 5.0449517E-13 alpha1 = -4.0583656E-18 beta0 = 6.2016506
+ aigbacc = 0.43 bigbacc = 0.054 cigbacc = 0.075
+ nigbacc = 1 aigbinv = 0.35 bigbinv = 0.03
+ cigbinv = 6E-3 eigbinv = 1.1 nigbinv = 3
+ aigc = 0.43 bigc = 0.054 cigc = 0.075
+ aigsd = 0.43 bigsd = 0.054 cigsd = 0.075
+ dlcig = 0 nigc = 1 poxedge = 1
+ pigcd = 1 ntox = 1 toxref = 4.23E-9
+ agidl = 0 bgidl = 2.3E9 cgidl = 0.5
+ egidl = 0.8 noia = 3E41 noib = 0
+ noic = 0 em = 4.1E7 af = 1
+ ef = 0.88 kf = 0 lintnoi = 0
+ tnoia = 2.5E7 tnoib = 0 ntnoi = 1
+ rnoia = 0.69 rnoib = 0.34 xpart = 0
+ cgso = {2E-11/sw_func_tox_lv_ratio} cgdo = {2E-11/sw_func_tox_lv_ratio} cgbo = {1E-13/sw_func_tox_lv_ratio}
+ ckappas = 0.6 cf = 0 clc = 7E-8
+ cle = 0.492 dlc = -1.2E-8 dwc = 0
+ vfbcv = -1 noff = 2.6123 voffcv = 0.112
+ acde = 0.44 moin = 8.7 cgsl = {0/sw_func_tox_lv_ratio}
+ cgdl = {0/sw_func_tox_lv_ratio} ijthsrev = 0.1 ijthsfwd = 0.1
+ xjbvs = 1 bvs = 12.69 jss = 2.1483E-5
+ jsws = 1.4472E-10 cjs = {7.682E-04*sw_func_psd_nw_cj} mjs = 0.3362
+ mjsws = 0.2659 cjsws = {9.160236799999998E-11*sw_func_psd_nw_cj} cjswgs = {2.39155046E-10*sw_func_psd_nw_cj}
+ mjswgs = 0.9274 pbs = 0.6587 pbsws = 0.7418
+ pbswgs = 1.4338 xrcrg1 = 12 xrcrg2 = 1
+ rbpb = 50 rbpd = 50 rbps = 50
+ rbdb = 50 rbsb = 50 gbmin = 1E-12
+ tnom = 30 ute = -0.312314378 lute = 7.163332394831999E-7
+ kt1 = -0.611336 lkt1 = 7.983207840000006E-8 kt1l = 0
+ kt2 = -0.055045 ua1 = 6.68269488E-10 lua1 = 1.111262531327999E-16
+ ub1 = -1.75362536E-19 lub1 = 2.136306417984E-25 uc1 = -9.961E-12
+ at = 2.99170974E5 lat = -0.1084917945456 prt = 0
+ njs = 1.3632 xtis = 5.2 tpb = 1.671E-3
+ tpbsw = 1.246E-3 tpbswg = 0 tcj = 1.2407E-3
+ tcjsw = 3.7357E-4 tcjswg = 2E-12 tvoff = 0
+ tvfbsdoff = 0 saref = 3E-6 sbref = 3E-6
+ wlod = 0 ku0 = 5.9E-8 kvsat = 0
+ kvth0 = 1.76E-8 tku0 = 0 llodku0 = 0
+ wlodku0 = 1 llodvth = 0 wlodvth = 1
+ lku0 = 0 wku0 = 0 pku0 = 0
+ lkvth0 = 0 wkvth0 = 7.3E-7 pkvth0 = 0
+ stk2 = 0 lodk2 = 1 steta0 = 0
+ lodeta0 = 1

.model plowvt_model.10 pmos
+ level = 54 lmin = 2E-6 lmax = 4E-6 wmin = 5E-6
+ wmax = 7E-6 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 4.23E-9
+ toxm = 4.23E-9 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 9.999999999999999E22 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {7.476E-9+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {2.8E-9-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = -7.916E-9 dwb = 0 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = -0.397075939860129 lvth0 = -3.109043406557387E-7
+ wvth0 = -1.767785764617417E-7 pvth0 = 1.594550234635303E-12 k1 = 0.64774
+ k2 = -0.024892036314955 lk2 = -9.051884911454258E-8 wk2 = -1.033409112670889E-7
+ pk2 = 4.362769332444949E-13 k3 = 3.39 k3b = 1
+ w0 = 1E-8 lpe0 = 0 lpeb = 0
+ vbm = -3 dvtp0 = 0 dvtp1 = 0
+ dvt0 = 2.4422 dvt1 = 0.16136 dvt2 = 0.026237
+ dvt0w = 0.5 dvt1w = 1.9281E6 dvt2w = -0.032
+ vfbsdoff = 0 u0 = 1.830227593137206E-3 lu0 = 4.015872579630434E-9
+ wu0 = 3.422796234320683E-9 pu0 = -1.985560055273532E-14 ua = -3.64520214549264E-9
+ lua = 2.91236073191612E-15 wua = 3.716534667427313E-15 pua = -1.569376410637883E-20
+ ub = 3.994770385390721E-18 lub = -4.290880125870933E-24 wub = -5.720035029411405E-24
+ pub = 2.374522682290815E-29 uc = 1.110001615482672E-10 luc = -7.867475725819692E-17
+ wuc = -3.466985627111336E-16 puc = 5.373883254985842E-22 ud = 0
+ up = 0 lp = 1 eu = 1.67
+ vsat = 2.387323757215936E5 lvsat = -0.459245657582333 wvsat = -0.573142811646179
+ pvsat = 2.289361646839496E-6 a0 = 3.513946250569836 la0 = -8.349591691208539E-6
+ wa0 = -8.739798589150373E-6 pa0 = 4.157883531844483E-11 ags = 0.691623993791211
+ lags = -1.225072978901032E-6 wags = -1.875740041833547E-6 pags = 7.956384720109313E-12
+ b0 = 0 b1 = 2.1073E-24 keta = -0.01258
+ a1 = 0 a2 = 0.46703705 rdsw = 484.7
+ rdswmin = 0 rdw = 0 rdwmin = 0
+ rsw = 0 rswmin = 0 prwb = 0.1
+ prwg = 0.052 wr = 1 voff = -0.1819
+ voffl = 0 minv = 0 nfactor = 2.5373
+ eta0 = 0.2 etab = -2.5E-4 dsub = 1
+ cit = -6.393105E-11 cdsc = 2.8125E-7 cdscb = 1E-4
+ cdscd = 1E-10 pclm = 0.030097 pdiblc1 = 0
+ pdiblc2 = 2.37520840416688E-3 lpdiblc2 = 9.814074073077412E-9 wpdiblc2 = -1.47481079982649E-8
+ ppdiblc2 = 2.511140955775421E-14 pdiblcb = -0.025 drout = 0.43496
+ pscbe1 = 8E8 pscbe2 = 8.6797E-9 pvag = 0
+ delta = 0.033465184523042 ldelta = -5.808546024870615E-8 wdelta = -9.62911479009843E-8
+ pdelta = 4.540303738597535E-13 fprout = 0 pdits = 0
+ pditsl = 0 pditsd = 0 lambda = 0
+ vtl = 0 lc = 5E-9 xn = 3
+ alpha0 = 5.0449517E-13 alpha1 = -4.0583656E-18 beta0 = 6.2016506
+ aigbacc = 0.43 bigbacc = 0.054 cigbacc = 0.075
+ nigbacc = 1 aigbinv = 0.35 bigbinv = 0.03
+ cigbinv = 6E-3 eigbinv = 1.1 nigbinv = 3
+ aigc = 0.43 bigc = 0.054 cigc = 0.075
+ aigsd = 0.43 bigsd = 0.054 cigsd = 0.075
+ dlcig = 0 nigc = 1 poxedge = 1
+ pigcd = 1 ntox = 1 toxref = 4.23E-9
+ agidl = 0 bgidl = 2.3E9 cgidl = 0.5
+ egidl = 0.8 noia = 3E41 noib = 0
+ noic = 0 em = 4.1E7 af = 1
+ ef = 0.88 kf = 0 lintnoi = 0
+ tnoia = 2.5E7 tnoib = 0 ntnoi = 1
+ rnoia = 0.69 rnoib = 0.34 xpart = 0
+ cgso = {2E-11/sw_func_tox_lv_ratio} cgdo = {2E-11/sw_func_tox_lv_ratio} cgbo = {1E-13/sw_func_tox_lv_ratio}
+ ckappas = 0.6 cf = 0 clc = 7E-8
+ cle = 0.492 dlc = -1.2E-8 dwc = 0
+ vfbcv = -1 noff = 2.6123 voffcv = 0.112
+ acde = 0.44 moin = 8.7 cgsl = {0/sw_func_tox_lv_ratio}
+ cgdl = {0/sw_func_tox_lv_ratio} ijthsrev = 0.1 ijthsfwd = 0.1
+ xjbvs = 1 bvs = 12.69 jss = 2.1483E-5
+ jsws = 1.4472E-10 cjs = {7.682E-04*sw_func_psd_nw_cj} mjs = 0.3362
+ mjsws = 0.2659 cjsws = {9.160236799999998E-11*sw_func_psd_nw_cj} cjswgs = {2.39155046E-10*sw_func_psd_nw_cj}
+ mjswgs = 0.9274 pbs = 0.6587 pbsws = 0.7418
+ pbswgs = 1.4338 xrcrg1 = 12 xrcrg2 = 1
+ rbpb = 50 rbpd = 50 rbps = 50
+ rbdb = 50 rbsb = 50 gbmin = 1E-12
+ tnom = 30 ute = -0.13298 kt1 = -0.59135
+ kt1l = 0 kt2 = -0.055045 ua1 = 6.9609E-10
+ ub1 = -2.44977619649816E-19 lub1 = 4.91701131929225E-25 wub1 = 6.13647542640076E-25
+ pub1 = -2.45115374432152E-30 uc1 = -9.961E-12 at = 5.81449301300352E5
+ lat = -1.236024345114126 wat = -1.420877490158829 pat = 5.675553046690426E-6
+ prt = 0 njs = 1.3632 xtis = 5.2
+ tpb = 1.671E-3 tpbsw = 1.246E-3 tpbswg = 0
+ tcj = 1.2407E-3 tcjsw = 3.7357E-4 tcjswg = 2E-12
+ tvoff = 0 tvfbsdoff = 0 saref = 3E-6
+ sbref = 3E-6 wlod = 0 ku0 = 5.9E-8
+ kvsat = 0 kvth0 = 1.76E-8 tku0 = 0
+ llodku0 = 0 wlodku0 = 1 llodvth = 0
+ wlodvth = 1 lku0 = 0 wku0 = 0
+ pku0 = 0 lkvth0 = 0 wkvth0 = 7.3E-7
+ pkvth0 = 0 stk2 = 0 lodk2 = 1
+ steta0 = 0 lodeta0 = 1

.model plowvt_model.11 pmos
+ level = 54 lmin = 1.5E-6 lmax = 2E-6 wmin = 5E-6
+ wmax = 7E-6 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 4.23E-9
+ toxm = 4.23E-9 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 9.999999999999999E22 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {7.476E-9+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {2.8E-9-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = -7.916E-9 dwb = 0 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = -0.629599509728205 lvth0 = 1.528406670891513E-7
+ wvth0 = 1.112083631123237E-6 pvth0 = -9.759565521721775E-13 k1 = 0.64774
+ k2 = -0.059219968731809 lk2 = -2.205522070236883E-8 wk2 = 8.168539499190612E-8
+ pk2 = 6.726046804155524E-14 k3 = 3.39 k3b = 1
+ w0 = 1E-8 lpe0 = 0 lpeb = 0
+ vbm = -3 dvtp0 = 0 dvtp1 = 0
+ dvt0 = 2.4422 dvt1 = 0.16136 dvt2 = 0.026237
+ dvt0w = 0.5 dvt1w = 1.9281E6 dvt2w = -0.032
+ vfbsdoff = 0 u0 = 5.342101449510924E-3 lu0 = -2.988208639521312E-9
+ wu0 = -1.527780319347085E-8 pu0 = 1.744087494605212E-14 ua = -4.901468211027183E-10
+ lua = -3.380081607047139E-15 wua = -1.218677007030082E-14 pua = 1.602378686254616E-20
+ ub = -8.162212032019188E-19 lub = 5.304161498418227E-24 wub = 1.849768064031692E-23
+ pub = -2.455458530879802E-29 uc = 5.303659098518401E-11 luc = 3.692778787281621E-17
+ wuc = -1.784603584031607E-16 puc = 2.018540508267631E-22 ud = 0
+ up = 0 lp = 1 eu = 1.67
+ vsat = -3.876929947617536E5 lvsat = 0.790097101309654 wvsat = 3.341933313578597
+ pvsat = -5.518866177308797E-6 a0 = -0.773096395755302 la0 = 2.004861626223164E-7
+ wa0 = 1.308767847755946E-5 pa0 = -1.953884943401262E-12 ags = 0.37104503872832
+ lags = -5.857103109236016E-7 wags = -1.423538356378182E-6 pags = 7.054513678637134E-12
+ b0 = 0 b1 = 2.1073E-24 keta = -0.01258
+ a1 = 0 a2 = 0.46703705 rdsw = 484.7
+ rdswmin = 0 rdw = 0 rdwmin = 0
+ rsw = 0 rswmin = 0 prwb = 0.1
+ prwg = 0.052 wr = 1 voff = -0.1819
+ voffl = 0 minv = 0 nfactor = 2.5373
+ eta0 = 0.2 etab = -2.5E-4 dsub = 1
+ cit = -6.393105E-11 cdsc = 2.8125E-7 cdscb = 1E-4
+ cdscd = 1E-10 pclm = 0.030097 pdiblc1 = 0
+ pdiblc2 = -6.755076593422732E-3 lpdiblc2 = 2.802351447227013E-8 wpdiblc2 = 2.428244614328272E-8
+ ppdiblc2 = -5.273112762214835E-14 pdiblcb = -0.025 drout = 0.43496
+ pscbe1 = 8E8 pscbe2 = 8.6797E-9 pvag = 0
+ delta = -6.396132487494385E-3 ldelta = 2.14139503971068E-8 wdelta = 1.632076225027269E-7
+ pdelta = -6.351397383340804E-14 fprout = 0 pdits = 0
+ pditsl = 0 pditsd = 0 lambda = 0
+ vtl = 0 lc = 5E-9 xn = 3
+ alpha0 = 5.0449517E-13 alpha1 = -4.0583656E-18 beta0 = 6.2016506
+ aigbacc = 0.43 bigbacc = 0.054 cigbacc = 0.075
+ nigbacc = 1 aigbinv = 0.35 bigbinv = 0.03
+ cigbinv = 6E-3 eigbinv = 1.1 nigbinv = 3
+ aigc = 0.43 bigc = 0.054 cigc = 0.075
+ aigsd = 0.43 bigsd = 0.054 cigsd = 0.075
+ dlcig = 0 nigc = 1 poxedge = 1
+ pigcd = 1 ntox = 1 toxref = 4.23E-9
+ agidl = 0 bgidl = 2.3E9 cgidl = 0.5
+ egidl = 0.8 noia = 3E41 noib = 0
+ noic = 0 em = 4.1E7 af = 1
+ ef = 0.88 kf = 0 lintnoi = 0
+ tnoia = 2.5E7 tnoib = 0 ntnoi = 1
+ rnoia = 0.69 rnoib = 0.34 xpart = 0
+ cgso = {2E-11/sw_func_tox_lv_ratio} cgdo = {2E-11/sw_func_tox_lv_ratio} cgbo = {1E-13/sw_func_tox_lv_ratio}
+ ckappas = 0.6 cf = 0 clc = 7E-8
+ cle = 0.492 dlc = -1.2E-8 dwc = 0
+ vfbcv = -1 noff = 2.6123 voffcv = 0.112
+ acde = 0.44 moin = 8.7 cgsl = {0/sw_func_tox_lv_ratio}
+ cgdl = {0/sw_func_tox_lv_ratio} ijthsrev = 0.1 ijthsfwd = 0.1
+ xjbvs = 1 bvs = 12.69 jss = 2.1483E-5
+ jsws = 1.4472E-10 cjs = {7.682E-04*sw_func_psd_nw_cj} mjs = 0.3362
+ mjsws = 0.2659 cjsws = {9.160236799999998E-11*sw_func_psd_nw_cj} cjswgs = {2.39155046E-10*sw_func_psd_nw_cj}
+ mjswgs = 0.9274 pbs = 0.6587 pbsws = 0.7418
+ pbswgs = 1.4338 xrcrg1 = 12 xrcrg2 = 1
+ rbpb = 50 rbpd = 50 rbps = 50
+ rbdb = 50 rbsb = 50 gbmin = 1E-12
+ tnom = 30 ute = -0.13298 kt1 = -0.814839671935999
+ lkt1 = 4.457278017091571E-7 wkt1 = 1.561086085977209E-6 pkt1 = -3.113430089872944E-12
+ kt1l = 0 kt2 = -0.206772138277351 lkt2 = 3.026046045803478E-7
+ wkt2 = 1.05982134376993E-6 pkt2 = -2.113707688014749E-12 ua1 = 8.464370986480642E-10
+ lua1 = -2.998522535436991E-16 wua1 = -3.236651818259424E-16 pua1 = 6.455178386336595E-22
+ ub1 = 3.893300659926387E-20 lub1 = -7.453022106194001E-26 wub1 = -2.454590170560303E-24
+ pub1 = 3.668139550885317E-30 uc1 = -9.961E-12 at = -8.460038989278721E5
+ lat = 1.610888317421044 wat = 7.347107366258367 pat = -1.181131595094803E-5
+ prt = 0 njs = 1.3632 xtis = 5.2
+ tpb = 1.671E-3 tpbsw = 1.246E-3 tpbswg = 0
+ tcj = 1.2407E-3 tcjsw = 3.7357E-4 tcjswg = 2E-12
+ tvoff = 0 tvfbsdoff = 0 saref = 3E-6
+ sbref = 3E-6 wlod = 0 ku0 = 5.9E-8
+ kvsat = 0 kvth0 = 1.76E-8 tku0 = 0
+ llodku0 = 0 wlodku0 = 1 llodvth = 0
+ wlodvth = 1 lku0 = 0 wku0 = 0
+ pku0 = 0 lkvth0 = 0 wkvth0 = 7.3E-7
+ pkvth0 = 0 stk2 = 0 lodk2 = 1
+ steta0 = 0 lodeta0 = 1

.model plowvt_model.12 pmos
+ level = 54 lmin = 1E-6 lmax = 1.5E-6 wmin = 5E-6
+ wmax = 7E-6 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 4.23E-9
+ toxm = 4.23E-9 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 9.999999999999999E22 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {7.476E-9+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {2.8E-9-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = -7.916E-9 dwb = 0 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = -0.499245780612538 lvth0 = -4.195994570130213E-8
+ wvth0 = 3.507328935842623E-7 pvth0 = 1.618059900060656E-13 k1 = 0.64774
+ k2 = -0.05528005725156 lk2 = -2.794302441845343E-8 wk2 = 2.917985900411621E-8
+ pk2 = 1.457247410217085E-13 k3 = 3.39 k3b = 1
+ w0 = 1E-8 lpe0 = 0 lpeb = 0
+ vbm = -3 dvtp0 = 0 dvtp1 = 0
+ dvt0 = 2.4422 dvt1 = 0.16136 dvt2 = 0.026237
+ dvt0w = 0.5 dvt1w = 1.9281E6 dvt2w = -0.032
+ vfbsdoff = 0 u0 = 1.765272969262423E-3 lu0 = 2.35700384136205E-9
+ wu0 = 1.843493199953384E-9 pu0 = -8.145190384281057E-15 ua = -3.222586688066563E-9
+ lua = 7.032765301436302E-16 wua = 4.852180920768445E-16 pua = -2.913232247311023E-21
+ ub = 3.124193357666559E-18 lub = -5.843940213436257E-25 wub = 1.171817403510353E-25
+ pub = 2.913232247310999E-30 uc = 1.04037491545088E-10 luc = -3.928795792390429E-17
+ wuc = -2.42138825961125E-16 puc = 2.97015152745385E-22 ud = 0
+ up = 0 lp = 1 eu = 1.67
+ vsat = 4.24755308978912E5 lvsat = -0.424025643800397 wvsat = -2.338099832005382
+ pvsat = 2.969375355451903E-6 a0 = -2.280614090763963 la0 = 2.453320606043259E-6
+ wa0 = 2.200409891475276E-5 pa0 = -1.527858364474292E-11 ags = -1.808012019458477
+ lags = 2.670672556830748E-6 wags = 1.24803421978759E-5 pags = -1.372344542164017E-11
+ b0 = 0 b1 = 2.1073E-24 keta = -0.01258
+ a1 = 0 a2 = 0.46703705 rdsw = 484.7
+ rdswmin = 0 rdw = 0 rdwmin = 0
+ rsw = 0 rswmin = 0 prwb = 0.1
+ prwg = 0.052 wr = 1 voff = -0.08083669331104
+ lvoff = -1.510290055159819E-7 wvoff = -5.03805434883187E-7 pvoff = 7.528868418894347E-13
+ voffl = 0 minv = 0 nfactor = 2.748456324628481
+ lnfactor = -3.155520115248027E-7 wnfactor = -1.052624413776562E-6 pnfactor = 1.573041923947695E-12
+ eta0 = 0.2 etab = -2.5E-4 dsub = 1
+ cit = -6.393105E-11 cdsc = 2.8125E-7 cdscb = 1E-4
+ cdscd = 1E-10 pclm = 0.030097 pdiblc1 = 0
+ pdiblc2 = 0.017390997582784 lpdiblc2 = -8.060378776653207E-9 wpdiblc2 = -1.173045881318862E-7
+ ppdiblc2 = 1.588565363986641E-13 pdiblcb = -0.025 drout = 0.43496
+ pscbe1 = 8E8 pscbe2 = 8.6797E-9 pvag = 0
+ delta = 5.502178719667187E-3 ldelta = 3.633114129124552E-9 wdelta = 3.306839407521171E-8
+ pdelta = 1.309660891286706E-13 fprout = 0 pdits = 0
+ pditsl = 0 pditsd = 0 lambda = 0
+ vtl = 0 lc = 5E-9 xn = 3
+ alpha0 = 5.0449517E-13 alpha1 = -4.0583656E-18 beta0 = 6.2016506
+ aigbacc = 0.43 bigbacc = 0.054 cigbacc = 0.075
+ nigbacc = 1 aigbinv = 0.35 bigbinv = 0.03
+ cigbinv = 6E-3 eigbinv = 1.1 nigbinv = 3
+ aigc = 0.43 bigc = 0.054 cigc = 0.075
+ aigsd = 0.43 bigsd = 0.054 cigsd = 0.075
+ dlcig = 0 nigc = 1 poxedge = 1
+ pigcd = 1 ntox = 1 toxref = 4.23E-9
+ agidl = 0 bgidl = 2.3E9 cgidl = 0.5
+ egidl = 0.8 noia = 3E41 noib = 0
+ noic = 0 em = 4.1E7 af = 1
+ ef = 0.88 kf = 0 lintnoi = 0
+ tnoia = 2.5E7 tnoib = 0 ntnoi = 1
+ rnoia = 0.69 rnoib = 0.34 xpart = 0
+ cgso = {2E-11/sw_func_tox_lv_ratio} cgdo = {2E-11/sw_func_tox_lv_ratio} cgbo = {1E-13/sw_func_tox_lv_ratio}
+ ckappas = 0.6 cf = 0 clc = 7E-8
+ cle = 0.492 dlc = -1.2E-8 dwc = 0
+ vfbcv = -1 noff = 2.6123 voffcv = 0.112
+ acde = 0.44 moin = 8.7 cgsl = {0/sw_func_tox_lv_ratio}
+ cgdl = {0/sw_func_tox_lv_ratio} ijthsrev = 0.1 ijthsfwd = 0.1
+ xjbvs = 1 bvs = 12.69 jss = 2.1483E-5
+ jsws = 1.4472E-10 cjs = {7.682E-04*sw_func_psd_nw_cj} mjs = 0.3362
+ mjsws = 0.2659 cjsws = {9.160236799999998E-11*sw_func_psd_nw_cj} cjswgs = {2.39155046E-10*sw_func_psd_nw_cj}
+ mjswgs = 0.9274 pbs = 0.6587 pbsws = 0.7418
+ pbswgs = 1.4338 xrcrg1 = 12 xrcrg2 = 1
+ rbpb = 50 rbpd = 50 rbps = 50
+ rbdb = 50 rbsb = 50 gbmin = 1E-12
+ tnom = 30 ute = 0.343024093284544 lute = -7.113405170044227E-7
+ wute = -2.003795224514778E-6 pute = 2.994471583514884E-12 kt1 = -0.625809597312001
+ lkt1 = 1.632412581910538E-7 wkt1 = -1.760539625870033E-7 pkt1 = -5.174480012985865E-13
+ kt1l = 0 kt2 = 0.058365917477351 lkt2 = -9.361770593947736E-8
+ wkt2 = -1.05982134376993E-6 pkt2 = 1.053886344244819E-12 ua1 = 5.166036478049278E-10
+ lua1 = 1.930508553962837E-16 wua1 = 1.010641115027484E-15 pua1 = -1.348469491384101E-21
+ ub1 = -9.418840950867203E-21 lub1 = -2.273220083024052E-27 wub1 = -7.583050875561352E-27
+ pub1 = 1.133211122843888E-32 uc1 = -9.961E-12 at = 9.371843411829124E5
+ lat = -1.053908188600512 wat = -5.118906295450762 pat = 6.817894865110094E-6
+ prt = 0 njs = 1.3632 xtis = 5.2
+ tpb = 1.671E-3 tpbsw = 1.246E-3 tpbswg = 0
+ tcj = 1.2407E-3 tcjsw = 3.7357E-4 tcjswg = 2E-12
+ tvoff = 0 tvfbsdoff = 0 saref = 3E-6
+ sbref = 3E-6 wlod = 0 ku0 = 5.9E-8
+ kvsat = 0 kvth0 = 1.76E-8 tku0 = 0
+ llodku0 = 0 wlodku0 = 1 llodvth = 0
+ wlodvth = 1 lku0 = 0 wku0 = 0
+ pku0 = 0 lkvth0 = 0 wkvth0 = 7.3E-7
+ pkvth0 = 0 stk2 = 0 lodk2 = 1
+ steta0 = 0 lodeta0 = 1

.model plowvt_model.13 pmos
+ level = 54 lmin = 5E-7 lmax = 1E-6 wmin = 5E-6
+ wmax = 7E-6 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 4.23E-9
+ toxm = 4.23E-9 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 9.999999999999999E22 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {7.476E-9+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {2.8E-9-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = -7.916E-9 dwb = 0 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = -0.570237732756627 lvth0 = 2.86344515107805E-8
+ wvth0 = 6.783908789977747E-7 pvth0 = -1.640171106891312E-13 k1 = 0.64774
+ k2 = -0.111795334189687 lk2 = 2.825576696881985E-8 wk2 = 3.365914916370652E-7
+ pk2 = -1.59965386468496E-13 k3 = 3.39 k3b = 1
+ w0 = 1E-8 lpe0 = 0 lpeb = 0
+ vbm = -3 dvtp0 = 0 dvtp1 = 0
+ dvt0 = 2.4422 dvt1 = 0.16136 dvt2 = 0.026237
+ dvt0w = 0.5 dvt1w = 1.9281E6 dvt2w = -0.032
+ vfbsdoff = 0 u0 = 5.222720487760016E-3 lu0 = -1.081081971031957E-9
+ wu0 = -1.382151051548685E-8 pu0 = 7.432089310352708E-15 ua = -1.77544594606848E-9
+ lua = -7.357602236992632E-16 wua = -7.085692859925136E-15 pua = 4.615281603359747E-21
+ ub = 1.488559255792641E-18 lub = 1.042080529559798E-24 wub = 9.335606788507807E-24
+ pub = -6.253569620576094E-30 uc = 3.651704314109443E-11 luc = 2.785437596902689E-17
+ wuc = 2.741172454401174E-16 puc = -2.163498846560105E-22 ud = 0
+ up = 0 lp = 1 eu = 1.67
+ vsat = 8.779420909536013E3 lvsat = -0.010379220704209 wvsat = 0.38064245614974
+ pvsat = 2.658580241104483E-7 a0 = 0.897442975297312 la0 = -7.069393404480723E-7
+ wa0 = 2.152536726907504E-6 pa0 = 4.461809794850398E-12 ags = 1.132073412325293
+ lags = -2.529483965350328E-7 wags = -1.247548937625242E-6 pags = -7.243047649783018E-14
+ b0 = -5.063575780573437E-7 lb0 = 5.035219756202227E-13 wb0 = 8.639894455979286E-12
+ pb0 = -8.591511047025801E-18 b1 = 2.1073E-24 keta = -0.01258
+ a1 = 0 a2 = 0.46703705 rdsw = 484.7
+ rdswmin = 0 rdw = 0 rdwmin = 0
+ rsw = 0 rswmin = 0 prwb = 0.1
+ prwg = 0.052 wr = 1 voff = -0.28296330668896
+ lvoff = 4.996569882702184E-8 wvoff = 5.038054348831869E-7 pvoff = -2.490814070062476E-13
+ voffl = 0 minv = 0 nfactor = 2.326143675371519
+ lnfactor = 1.043956868963212E-7 wnfactor = 1.052624413776562E-6 pnfactor = -5.204175101711322E-13
+ eta0 = 0.2 etab = -2.5E-4 dsub = 1
+ cit = -6.393105E-11 cdsc = 2.8125E-7 cdscb = 1E-4
+ cdscd = 1E-10 pclm = 0.030097 pdiblc1 = 0
+ pdiblc2 = -0.04153656098953 lpdiblc2 = 5.053718546765543E-8 wpdiblc2 = 1.312436049064333E-7
+ ppdiblc2 = -8.829978675864084E-14 pdiblcb = -0.025 drout = 0.43496
+ pscbe1 = 8E8 pscbe2 = 8.6797E-9 pvag = 0
+ delta = 4.10625690999041E-3 ldelta = 5.021218776667141E-9 wdelta = 1.205800832484734E-7
+ pdelta = 4.394446541477919E-14 fprout = 0 pdits = 0
+ pditsl = 0 pditsd = 0 lambda = 0
+ vtl = 0 lc = 5E-9 xn = 3
+ alpha0 = 5.0449517E-13 alpha1 = -4.0583656E-18 beta0 = 6.2016506
+ aigbacc = 0.43 bigbacc = 0.054 cigbacc = 0.075
+ nigbacc = 1 aigbinv = 0.35 bigbinv = 0.03
+ cigbinv = 6E-3 eigbinv = 1.1 nigbinv = 3
+ aigc = 0.43 bigc = 0.054 cigc = 0.075
+ aigsd = 0.43 bigsd = 0.054 cigsd = 0.075
+ dlcig = 0 nigc = 1 poxedge = 1
+ pigcd = 1 ntox = 1 toxref = 4.23E-9
+ agidl = 0 bgidl = 2.3E9 cgidl = 0.5
+ egidl = 0.8 noia = 3E41 noib = 0
+ noic = 0 em = 4.1E7 af = 1
+ ef = 0.88 kf = 0 lintnoi = 0
+ tnoia = 2.5E7 tnoib = 0 ntnoi = 1
+ rnoia = 0.69 rnoib = 0.34 xpart = 0
+ cgso = {2E-11/sw_func_tox_lv_ratio} cgdo = {2E-11/sw_func_tox_lv_ratio} cgbo = {1E-13/sw_func_tox_lv_ratio}
+ ckappas = 0.6 cf = 0 clc = 7E-8
+ cle = 0.492 dlc = -1.2E-8 dwc = 0
+ vfbcv = -1 noff = 2.6123 voffcv = 0.112
+ acde = 0.44 moin = 8.7 cgsl = {0/sw_func_tox_lv_ratio}
+ cgdl = {0/sw_func_tox_lv_ratio} ijthsrev = 0.1 ijthsfwd = 0.1
+ xjbvs = 1 bvs = 12.69 jss = 2.1483E-5
+ jsws = 1.4472E-10 cjs = {7.682E-04*sw_func_psd_nw_cj} mjs = 0.3362
+ mjsws = 0.2659 cjsws = {9.160236799999998E-11*sw_func_psd_nw_cj} cjswgs = {2.39155046E-10*sw_func_psd_nw_cj}
+ mjswgs = 0.9274 pbs = 0.6587 pbsws = 0.7418
+ pbswgs = 1.4338 xrcrg1 = 12 xrcrg2 = 1
+ rbpb = 50 rbpd = 50 rbps = 50
+ rbdb = 50 rbsb = 50 gbmin = 1E-12
+ tnom = 30 ute = -0.346457693284544 lute = -2.571982844012144E-8
+ wute = 2.003795224514778E-6 pute = -9.90676359000106E-13 kt1 = -0.308821883613184
+ lkt1 = -1.519713243110499E-7 wkt1 = -1.276230774511433E-6 pkt1 = 5.76567820479067E-13
+ kt1l = 0 kt2 = -0.0157696432 lkt2 = -1.989730440192E-8
+ ua1 = 5.27212165547008E-10 lua1 = 1.825017453535592E-16 wua1 = -6.869759332015413E-16
+ pua1 = 3.39640901374842E-22 ub1 = 5.692301049508672E-19 lub1 = -5.776817318877087E-25
+ wub1 = 7.58305087556135E-27 pub1 = -3.749060352877532E-33 uc1 = -2.284941472E-11
+ luc1 = 1.2816239597568E-17 at = -3.02615596256448E5 lat = 0.178948869189188
+ wat = 3.455308889827711 pat = -1.70830471513082E-6 prt = 0
+ njs = 1.3632 xtis = 5.2 tpb = 1.671E-3
+ tpbsw = 1.246E-3 tpbswg = 0 tcj = 1.2407E-3
+ tcjsw = 3.7357E-4 tcjswg = 2E-12 tvoff = 0
+ tvfbsdoff = 0 saref = 2.74E-6 sbref = 2.74E-6
+ wlod = 0 ku0 = 5.9E-8 kvsat = 0
+ kvth0 = 1.76E-8 tku0 = 0 llodku0 = 0
+ wlodku0 = 1 llodvth = 0 wlodvth = 1
+ lku0 = 0 wku0 = 0 pku0 = 0
+ lkvth0 = 0 wkvth0 = 7.3E-7 pkvth0 = 0
+ stk2 = 0 lodk2 = 1 steta0 = 0
+ lodeta0 = 1

.model plowvt_model.14 pmos
+ level = 54 lmin = 3.5E-7 lmax = 5E-7 wmin = 5E-6
+ wmax = 7E-6 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 4.23E-9
+ toxm = 4.23E-9 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 9.999999999999999E22 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {7.476E-9+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {2.8E-9-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = -7.916E-9 dwb = 0 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = -0.564898394654784 lvth0 = 2.59946827532293E-8
+ wvth0 = 5.983191132855544E-7 pvth0 = -1.244296297210094E-13 k1 = 0.64774
+ k2 = -0.060038015441581 lk2 = 2.666948579756257E-9 wk2 = -4.331882962380421E-8
+ pk2 = 2.786227636287781E-14 k3 = 3.39 k3b = 1
+ w0 = 1E-8 lpe0 = 0 lpeb = 0
+ vbm = -3 dvtp0 = 0 dvtp1 = 0
+ dvt0 = 2.4422 dvt1 = 0.16136 dvt2 = 0.026237
+ dvt0w = 0.5 dvt1w = 1.9281E6 dvt2w = -0.032
+ vfbsdoff = 0 u0 = 1.348473446949025E-3 lu0 = 8.343457659449974E-10
+ wu0 = 7.377824464950646E-9 pu0 = -3.048861903975588E-15 ua = -4.135503596236799E-9
+ lua = 4.310522785439536E-16 wua = 7.414100356085063E-15 pua = -2.553416162635696E-21
+ ub = 4.593542837491201E-18 lub = -4.930233532319697E-25 wub = -1.092030416225224E-23
+ pub = 3.76095275347967E-30 uc = 1.610911659865599E-10 luc = -3.373507036577124E-17
+ wuc = -5.388421234027765E-16 puc = 1.855772272999162E-22 ud = 0
+ up = 0 lp = 1 eu = 1.67
+ vsat = -2.612834642092352E5 lvsat = 0.123139869698512 wvsat = 2.930638358283918
+ pvsat = -9.94859949904689E-7 a0 = -4.050956889740545 la0 = 1.739549552826643E-6
+ wa0 = 3.684015968422313E-5 pa0 = -1.268775099524644E-11 ags = 1.09346676605344
+ lags = -2.338612706182289E-7 wags = -4.766280793912052E-6 pags = 1.667230553250368E-12
+ b0 = 1.68785859352448E-6 lb0 = -5.81298499609831E-13 wb0 = -2.879964818659762E-11
+ pb0 = 9.91859883546422E-18 b1 = 2.1073E-24 keta = -0.01258
+ a1 = 0 a2 = 0.46703705 rdsw = 484.7
+ rdswmin = 0 rdw = 0 rdwmin = 0
+ rsw = 0 rswmin = 0 prwb = 0.1
+ prwg = 0.052 wr = 1 voff = -0.1819
+ voffl = 0 minv = 0 nfactor = 2.5373
+ eta0 = 0.2 etab = -2.5E-4 dsub = 1
+ cit = -6.393105E-11 cdsc = 2.8125E-7 cdscb = 1E-4
+ cdscd = 1E-10 pclm = 0.030097 pdiblc1 = 0
+ pdiblc2 = -0.15762177437456 lpdiblc2 = 1.079297149652145E-7 wpdiblc2 = 4.829025089059355E-7
+ ppdiblc2 = -2.621599488959947E-13 pdiblcb = -0.025 drout = 0.43496
+ pscbe1 = 8E8 pscbe2 = 8.6797E-9 pvag = 0
+ delta = 1.42776893945605E-3 ldelta = 6.345463229299331E-9 wdelta = 1.639338172417584E-7
+ pdelta = 2.251037932849907E-14 fprout = 0 pdits = 0
+ pditsl = 0 pditsd = 0 lambda = 0
+ vtl = 0 lc = 5E-9 xn = 3
+ alpha0 = 5.0449517E-13 alpha1 = -4.0583656E-18 beta0 = 6.2016506
+ aigbacc = 0.43 bigbacc = 0.054 cigbacc = 0.075
+ nigbacc = 1 aigbinv = 0.35 bigbinv = 0.03
+ cigbinv = 6E-3 eigbinv = 1.1 nigbinv = 3
+ aigc = 0.43 bigc = 0.054 cigc = 0.075
+ aigsd = 0.43 bigsd = 0.054 cigsd = 0.075
+ dlcig = 0 nigc = 1 poxedge = 1
+ pigcd = 1 ntox = 1 toxref = 4.23E-9
+ agidl = 0 bgidl = 2.3E9 cgidl = 0.5
+ egidl = 0.8 noia = 3E41 noib = 0
+ noic = 0 em = 4.1E7 af = 1
+ ef = 0.88 kf = 0 lintnoi = 0
+ tnoia = 2.5E7 tnoib = 0 ntnoi = 1
+ rnoia = 0.69 rnoib = 0.34 xpart = 0
+ cgso = {2E-11/sw_func_tox_lv_ratio} cgdo = {2E-11/sw_func_tox_lv_ratio} cgbo = {1E-13/sw_func_tox_lv_ratio}
+ ckappas = 0.6 cf = 0 clc = 7E-8
+ cle = 0.492 dlc = -1.2E-8 dwc = 0
+ vfbcv = -1 noff = 2.6123 voffcv = 0.112
+ acde = 0.44 moin = 8.7 cgsl = {0/sw_func_tox_lv_ratio}
+ cgdl = {0/sw_func_tox_lv_ratio} ijthsrev = 0.1 ijthsfwd = 0.1
+ xjbvs = 1 bvs = 12.69 jss = 2.1483E-5
+ jsws = 1.4472E-10 cjs = {7.682E-04*sw_func_psd_nw_cj} mjs = 0.3362
+ mjsws = 0.2659 cjsws = {9.160236799999998E-11*sw_func_psd_nw_cj} cjswgs = {2.39155046E-10*sw_func_psd_nw_cj}
+ mjswgs = 0.9274 pbs = 0.6587 pbsws = 0.7418
+ pbswgs = 1.4338 xrcrg1 = 12 xrcrg2 = 1
+ rbpb = 50 rbpd = 50 rbps = 50
+ rbdb = 50 rbsb = 50 gbmin = 1E-12
+ tnom = 30 ute = -0.39848 kt1 = -0.60299893046272
+ lkt1 = -6.530192348639202E-9 wkt1 = -3.626711629292382E-7 pkt1 = 1.249039485128296E-13
+ kt1l = 0 kt2 = -0.056015 ua1 = 8.9635E-10
+ ub1 = -5.9922E-19 uc1 = 3.0734E-12 at = 1.37677816E5
+ lat = -0.0387321938304 prt = 0 njs = 1.3632
+ xtis = 5.2 tpb = 1.671E-3 tpbsw = 1.246E-3
+ tpbswg = 0 tcj = 1.2407E-3 tcjsw = 3.7357E-4
+ tcjswg = 2E-12 tvoff = 0 tvfbsdoff = 0
+ saref = 1.74E-6 sbref = 1.74E-6 wlod = 0
+ ku0 = 5.9E-8 kvsat = 0 kvth0 = 1.76E-8
+ tku0 = 0 llodku0 = 0 wlodku0 = 1
+ llodvth = 0 wlodvth = 1 lku0 = 0
+ wku0 = 0 pku0 = 0 lkvth0 = 0
+ wkvth0 = 7.3E-7 pkvth0 = 0 stk2 = 0
+ lodk2 = 1 steta0 = 0 lodeta0 = 1

.model plowvt_model.15 pmos
+ level = 54 lmin = 8E-6 lmax = 2.02E-5 wmin = 3E-6
+ wmax = 5E-6 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 4.23E-9
+ toxm = 4.23E-9 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 9.999999999999999E22 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {7.476E-9+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {2.8E-9-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = -7.916E-9 dwb = 0 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = -0.4449641246552 wvth0 = 3.042935440415529E-8
+ k1 = 0.64774 k2 = -0.0442445335312 wk2 = -7.895650372558493E-9
+ k3 = 3.39 k3b = 1 w0 = 1E-8
+ lpe0 = 0 lpeb = 0 vbm = -3
+ dvtp0 = 0 dvtp1 = 0 dvt0 = 2.4422
+ dvt1 = 0.16136 dvt2 = 0.026237 dvt0w = 0.5
+ dvt1w = 1.9281E6 dvt2w = -0.032 vfbsdoff = 0
+ u0 = 2.148846436628E-3 wu0 = 1.770442605636462E-9 ua = -3.1079524E-9
+ wua = 7.440303781152008E-16 ub = 3.07007668E-18 wub = -5.208212646806403E-25
+ uc = 3.055610253599999E-11 wuc = 9.066754187711833E-17 ud = 0
+ up = 0 lp = 1 eu = 1.67
+ vsat = 1.2376E5 a0 = 1.766947498856 wa0 = -6.319794031710512E-8
+ ags = 0.373610259156 wags = -4.701527959309923E-8 b0 = 0
+ b1 = 2.1073E-24 keta = -0.01258 a1 = 0
+ a2 = 0.46703705 rdsw = 484.7 rdswmin = 0
+ rdw = 0 rdwmin = 0 rsw = 0
+ rswmin = 0 prwb = 0.1 prwg = 0.052
+ wr = 1 voff = -0.1819 voffl = 0
+ minv = 0 nfactor = 2.5373 eta0 = 0.2
+ etab = -2.5E-4 dsub = 1 cit = -6.393105E-11
+ cdsc = 2.8125E-7 cdscb = 1E-4 cdscd = 1E-10
+ pclm = 0.030097 pdiblc1 = 0 pdiblc2 = 7.438602707999997E-4
+ wpdiblc2 = 4.488735271169004E-9 pdiblcb = -0.025 drout = 0.43496
+ pscbe1 = 8E8 pscbe2 = 8.6797E-9 pvag = 0
+ delta = 0.013271681292 wdelta = 2.2075381318678E-8 fprout = 0
+ pdits = 0 pditsl = 0 pditsd = 0
+ lambda = 0 vtl = 0 lc = 5E-9
+ xn = 3 alpha0 = 5.0449517E-13 alpha1 = -4.0583656E-18
+ beta0 = 6.2016506 aigbacc = 0.43 bigbacc = 0.054
+ cigbacc = 0.075 nigbacc = 1 aigbinv = 0.35
+ bigbinv = 0.03 cigbinv = 6E-3 eigbinv = 1.1
+ nigbinv = 3 aigc = 0.43 bigc = 0.054
+ cigc = 0.075 aigsd = 0.43 bigsd = 0.054
+ cigsd = 0.075 dlcig = 0 nigc = 1
+ poxedge = 1 pigcd = 1 ntox = 1
+ toxref = 4.23E-9 agidl = 0 bgidl = 2.3E9
+ cgidl = 0.5 egidl = 0.8 noia = 3E41
+ noib = 0 noic = 0 em = 4.1E7
+ af = 1 ef = 0.88 kf = 0
+ lintnoi = 0 tnoia = 2.5E7 tnoib = 0
+ ntnoi = 1 rnoia = 0.69 rnoib = 0.34
+ xpart = 0 cgso = {2E-11/sw_func_tox_lv_ratio} cgdo = {2E-11/sw_func_tox_lv_ratio}
+ cgbo = {1E-13/sw_func_tox_lv_ratio} ckappas = 0.6 cf = 0
+ clc = 7E-8 cle = 0.492 dlc = -1.2E-8
+ dwc = 0 vfbcv = -1 noff = 2.6123
+ voffcv = 0.112 acde = 0.44 moin = 8.7
+ cgsl = {0/sw_func_tox_lv_ratio} cgdl = {0/sw_func_tox_lv_ratio} ijthsrev = 0.1
+ ijthsfwd = 0.1 xjbvs = 1 bvs = 12.69
+ jss = 2.1483E-5 jsws = 1.4472E-10 cjs = {7.682E-04*sw_func_psd_nw_cj}
+ mjs = 0.3362 mjsws = 0.2659 cjsws = {9.160236799999998E-11*sw_func_psd_nw_cj}
+ cjswgs = {2.39155046E-10*sw_func_psd_nw_cj} mjswgs = 0.9274 pbs = 0.6587
+ pbsws = 0.7418 pbswgs = 1.4338 xrcrg1 = 12
+ xrcrg2 = 1 rbpb = 50 rbpd = 50
+ rbps = 50 rbdb = 50 rbsb = 50
+ gbmin = 1E-12 tnom = 30 ute = -0.11966614304
+ wute = -5.136785730507344E-7 kt1 = -0.60135 kt1l = 0
+ kt2 = -0.055045 ua1 = 6.8217E-10 ub1 = -1.4641613924E-19
+ wub1 = -1.108605263391646E-26 uc1 = -9.961E-12 at = 2.8986861864E5
+ wat = -0.021279268814095 prt = 0 njs = 1.3632
+ xtis = 5.2 tpb = 1.671E-3 tpbsw = 1.246E-3
+ tpbswg = 0 tcj = 1.2407E-3 tcjsw = 3.7357E-4
+ tcjswg = 2E-12 tvoff = 0 tvfbsdoff = 0
+ saref = 3E-6 sbref = 3E-6 wlod = 0
+ ku0 = 5.9E-8 kvsat = 0 kvth0 = 1.76E-8
+ tku0 = 0 llodku0 = 0 wlodku0 = 1
+ llodvth = 0 wlodvth = 1 lku0 = 0
+ wku0 = 0 pku0 = 0 lkvth0 = 0
+ wkvth0 = 7.3E-7 pkvth0 = 0 stk2 = 0
+ lodk2 = 1 steta0 = 0 lodeta0 = 1

.model plowvt_model.16 pmos
+ level = 54 lmin = 4E-6 lmax = 8E-6 wmin = 3E-6
+ wmax = 5E-6 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 4.23E-9
+ toxm = 4.23E-9 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 9.999999999999999E22 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {7.476E-9+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {2.8E-9-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = -7.916E-9 dwb = 0 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = -0.43876104251648 lvth0 = -4.958991984978157E-8
+ wvth0 = -4.31354462836702E-8 pvth0 = 5.88106442618752E-13 k1 = 0.64774
+ k2 = -0.036874254225428 lk2 = -5.892096088206422E-8 wk2 = -4.19223054961831E-8
+ pk2 = 2.720226917203045E-13 k3 = 3.39 k3b = 1
+ w0 = 1E-8 lpe0 = 0 lpeb = 0
+ vbm = -3 dvtp0 = 0 dvtp1 = 0
+ dvt0 = 2.4422 dvt1 = 0.16136 dvt2 = 0.026237
+ dvt0w = 0.5 dvt1w = 1.9281E6 dvt2w = -0.032
+ vfbsdoff = 0 u0 = 1.895206272629284E-3 lu0 = 2.027700927071333E-9
+ wu0 = 2.929987975828501E-9 pu0 = -9.269869507463237E-15 ua = -3.152665433992E-9
+ lua = 3.574538789456462E-16 wua = 9.669269987909532E-16 pua = -1.781924744330235E-21
+ ub = 3.07007668E-18 wub = -5.208212646806403E-25 uc = 3.055610253599999E-11
+ wuc = 9.066754187711833E-17 ud = 0 up = 0
+ lp = 1 eu = 1.67 vsat = 1.2376E5
+ a0 = 1.823456538575397 la0 = -4.517558671327448E-7 wa0 = -3.660550087166045E-7
+ pa0 = 2.421160547612958E-12 ags = 0.320883034976097 lags = 4.215225209838124E-7
+ wags = -3.431560363633635E-9 pags = -3.484256850080397E-13 b0 = 0
+ b1 = 2.1073E-24 keta = -0.01258 a1 = 0
+ a2 = 0.46703705 rdsw = 484.7 rdswmin = 0
+ rdw = 0 rdwmin = 0 rsw = 0
+ rswmin = 0 prwb = 0.1 prwg = 0.052
+ wr = 1 voff = -0.1819 voffl = 0
+ minv = 0 nfactor = 2.5373 eta0 = 0.2
+ etab = -2.5E-4 dsub = 1 cit = -6.393105E-11
+ cdsc = 2.8125E-7 cdscb = 1E-4 cdscd = 1E-10
+ pclm = 0.030097 pdiblc1 = 0 pdiblc2 = -1.49752052162528E-3
+ lpdiblc2 = 1.791849460696466E-8 wpdiblc2 = 8.242314363348664E-9 ppdiblc2 = -3.000761269452108E-14
+ pdiblcb = -0.025 drout = 0.43496 pscbe1 = 8E8
+ pscbe2 = 8.6797E-9 pvag = 0 delta = 0.011818421028752
+ ldelta = 1.161794384850977E-8 wdelta = 5.878226882906701E-9 pdelta = 1.294865314213301E-13
+ fprout = 0 pdits = 0 pditsl = 0
+ pditsd = 0 lambda = 0 vtl = 0
+ lc = 5E-9 xn = 3 alpha0 = 5.0449517E-13
+ alpha1 = -4.0583656E-18 beta0 = 6.2016506 aigbacc = 0.43
+ bigbacc = 0.054 cigbacc = 0.075 nigbacc = 1
+ aigbinv = 0.35 bigbinv = 0.03 cigbinv = 6E-3
+ eigbinv = 1.1 nigbinv = 3 aigc = 0.43
+ bigc = 0.054 cigc = 0.075 aigsd = 0.43
+ bigsd = 0.054 cigsd = 0.075 dlcig = 0
+ nigc = 1 poxedge = 1 pigcd = 1
+ ntox = 1 toxref = 4.23E-9 agidl = 0
+ bgidl = 2.3E9 cgidl = 0.5 egidl = 0.8
+ noia = 3E41 noib = 0 noic = 0
+ em = 4.1E7 af = 1 ef = 0.88
+ kf = 0 lintnoi = 0 tnoia = 2.5E7
+ tnoib = 0 ntnoi = 1 rnoia = 0.69
+ rnoib = 0.34 xpart = 0 cgso = {2E-11/sw_func_tox_lv_ratio}
+ cgdo = {2E-11/sw_func_tox_lv_ratio} cgbo = {1E-13/sw_func_tox_lv_ratio} ckappas = 0.6
+ cf = 0 clc = 7E-8 cle = 0.492
+ dlc = -1.2E-8 dwc = 0 vfbcv = -1
+ noff = 2.6123 voffcv = 0.112 acde = 0.44
+ moin = 8.7 cgsl = {0/sw_func_tox_lv_ratio} cgdl = {0/sw_func_tox_lv_ratio}
+ ijthsrev = 0.1 ijthsfwd = 0.1 xjbvs = 1
+ bvs = 12.69 jss = 2.1483E-5 jsws = 1.4472E-10
+ cjs = {7.682E-04*sw_func_psd_nw_cj} mjs = 0.3362 mjsws = 0.2659
+ cjsws = {9.160236799999998E-11*sw_func_psd_nw_cj} cjswgs = {2.39155046E-10*sw_func_psd_nw_cj} mjswgs = 0.9274
+ pbs = 0.6587 pbsws = 0.7418 pbswgs = 1.4338
+ xrcrg1 = 12 xrcrg2 = 1 rbpb = 50
+ rbpd = 50 rbps = 50 rbdb = 50
+ rbsb = 50 gbmin = 1E-12 tnom = 30
+ ute = -0.106370925479744 lute = -1.062872872637111E-7 wute = -1.026637996099198E-6
+ pute = 4.100802811618635E-12 kt1 = -0.611336 lkt1 = 7.983207840000006E-8
+ kt1l = 0 kt2 = -0.055045 ua1 = 6.68269488E-10
+ lua1 = 1.111262531327999E-16 ub1 = -1.70917927885064E-19 lub1 = 1.958770991440997E-25
+ wub1 = -2.215658479414543E-26 pub1 = 8.850226230173451E-32 uc1 = -9.961E-12
+ at = 3.07702235213904E5 lat = -0.142569064338418 wat = -0.04252874665185
+ pat = 1.698768256261485E-7 prt = 0 njs = 1.3632
+ xtis = 5.2 tpb = 1.671E-3 tpbsw = 1.246E-3
+ tpbswg = 0 tcj = 1.2407E-3 tcjsw = 3.7357E-4
+ tcjswg = 2E-12 tvoff = 0 tvfbsdoff = 0
+ saref = 3E-6 sbref = 3E-6 wlod = 0
+ ku0 = 5.9E-8 kvsat = 0 kvth0 = 1.76E-8
+ tku0 = 0 llodku0 = 0 wlodku0 = 1
+ llodvth = 0 wlodvth = 1 lku0 = 0
+ wku0 = 0 pku0 = 0 lkvth0 = 0
+ wkvth0 = 7.3E-7 pkvth0 = 0 stk2 = 0
+ lodk2 = 1 steta0 = 0 lodeta0 = 1

.model plowvt_model.17 pmos
+ level = 54 lmin = 2E-6 lmax = 4E-6 wmin = 3E-6
+ wmax = 5E-6 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 4.23E-9
+ toxm = 4.23E-9 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 9.999999999999999E22 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {7.476E-9+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {2.8E-9-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = -7.916E-9 dwb = 0 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = -0.447214693259157 lvth0 = -1.58226573232331E-8
+ wvth0 = 7.316551589257391E-8 pvth0 = 1.235538793019626E-13 k1 = 0.64774
+ k2 = -0.055667912471535 lk2 = 1.614842761618721E-8 wk2 = 5.007830861551849E-8
+ pk2 = -9.546456128747625E-14 k3 = 3.39 k3b = 1
+ w0 = 1E-8 lpe0 = 0 lpeb = 0
+ vbm = -3 dvtp0 = 0 dvtp1 = 0
+ dvt0 = 2.4422 dvt1 = 0.16136 dvt2 = 0.026237
+ dvt0w = 0.5 dvt1w = 1.9281E6 dvt2w = -0.032
+ vfbsdoff = 0 u0 = 2.375100636894328E-3 lu0 = 1.108108784510421E-10
+ wu0 = 7.065779572853304E-10 pu0 = -3.886805293943961E-16 ua = -2.91603241997824E-9
+ lua = -5.877530322309179E-16 wua = 8.158858559120537E-17 pua = 1.754471013354837E-21
+ ub = 2.775291050969919E-18 lub = 1.177491716597754E-24 wub = 3.591279876843443E-25
+ pub = -3.514869293646694E-30 uc = -2.128076762500812E-12 luc = 1.305536857899316E-16
+ wuc = 2.17251135423484E-16 puc = -5.056255060616031E-22 ud = 0
+ up = 0 lp = 1 eu = 1.67
+ vsat = 1.2376E5 a0 = 1.38801217034764 la0 = 1.287583117316204E-6
+ wa0 = 1.858084845593125E-6 pa0 = -6.462943686441824E-12 ags = 0.217959757183416
+ lags = 8.326392617988995E-7 wags = 4.854989135396709E-7 pags = -2.301409569967399E-12
+ b0 = 0 b1 = 2.1073E-24 keta = -0.01258
+ a1 = 0 a2 = 0.46703705 rdsw = 484.7
+ rdswmin = 0 rdw = 0 rdwmin = 0
+ rsw = 0 rswmin = 0 prwb = 0.1
+ prwg = 0.052 wr = 1 voff = -0.1819
+ voffl = 0 minv = 0 nfactor = 2.5373
+ eta0 = 0.2 etab = -2.5E-4 dsub = 1
+ cit = -6.393105E-11 cdsc = 2.8125E-7 cdscb = 1E-4
+ cdscd = 1E-10 pclm = 0.030097 pdiblc1 = 0
+ pdiblc2 = -1.46730055309568E-3 lpdiblc2 = 1.779778396467002E-8 wpdiblc2 = 4.406983594118915E-9
+ ppdiblc2 = -1.468776746990976E-14 pdiblcb = -0.025 drout = 0.43496
+ pscbe1 = 8E8 pscbe2 = 8.6797E-9 pvag = 0
+ delta = 0.012660174637381 ldelta = 8.25564323420298E-9 wdelta = 7.422825019509374E-9
+ pdelta = 1.233167886244843E-13 fprout = 0 pdits = 0
+ pditsl = 0 pditsd = 0 lambda = 0
+ vtl = 0 lc = 5E-9 xn = 3
+ alpha0 = 5.0449517E-13 alpha1 = -4.0583656E-18 beta0 = 6.2016506
+ aigbacc = 0.43 bigbacc = 0.054 cigbacc = 0.075
+ nigbacc = 1 aigbinv = 0.35 bigbinv = 0.03
+ cigbinv = 6E-3 eigbinv = 1.1 nigbinv = 3
+ aigc = 0.43 bigc = 0.054 cigc = 0.075
+ aigsd = 0.43 bigsd = 0.054 cigsd = 0.075
+ dlcig = 0 nigc = 1 poxedge = 1
+ pigcd = 1 ntox = 1 toxref = 4.23E-9
+ agidl = 0 bgidl = 2.3E9 cgidl = 0.5
+ egidl = 0.8 noia = 3E41 noib = 0
+ noic = 0 em = 4.1E7 af = 1
+ ef = 0.88 kf = 0 lintnoi = 0
+ tnoia = 2.5E7 tnoib = 0 ntnoi = 1
+ rnoia = 0.69 rnoib = 0.34 xpart = 0
+ cgso = {2E-11/sw_func_tox_lv_ratio} cgdo = {2E-11/sw_func_tox_lv_ratio} cgbo = {1E-13/sw_func_tox_lv_ratio}
+ ckappas = 0.6 cf = 0 clc = 7E-8
+ cle = 0.492 dlc = -1.2E-8 dwc = 0
+ vfbcv = -1 noff = 2.6123 voffcv = 0.112
+ acde = 0.44 moin = 8.7 cgsl = {0/sw_func_tox_lv_ratio}
+ cgdl = {0/sw_func_tox_lv_ratio} ijthsrev = 0.1 ijthsfwd = 0.1
+ xjbvs = 1 bvs = 12.69 jss = 2.1483E-5
+ jsws = 1.4472E-10 cjs = {7.682E-04*sw_func_psd_nw_cj} mjs = 0.3362
+ mjsws = 0.2659 cjsws = {9.160236799999998E-11*sw_func_psd_nw_cj} cjswgs = {2.39155046E-10*sw_func_psd_nw_cj}
+ mjswgs = 0.9274 pbs = 0.6587 pbsws = 0.7418
+ pbswgs = 1.4338 xrcrg1 = 12 xrcrg2 = 1
+ rbpb = 50 rbpd = 50 rbps = 50
+ rbdb = 50 rbsb = 50 gbmin = 1E-12
+ tnom = 30 ute = -0.13298 kt1 = -0.59135
+ kt1l = 0 kt2 = -0.055045 ua1 = 6.9609E-10
+ ub1 = -1.2188E-19 uc1 = -9.961E-12 at = 2.85363053149296E5
+ lat = -0.053337435499548 wat = 0.055126669014096 pat = -2.201979667099062E-7
+ prt = 0 njs = 1.3632 xtis = 5.2
+ tpb = 1.671E-3 tpbsw = 1.246E-3 tpbswg = 0
+ tcj = 1.2407E-3 tcjsw = 3.7357E-4 tcjswg = 2E-12
+ tvoff = 0 tvfbsdoff = 0 saref = 3E-6
+ sbref = 3E-6 wlod = 0 ku0 = 5.9E-8
+ kvsat = 0 kvth0 = 1.76E-8 tku0 = 0
+ llodku0 = 0 wlodku0 = 1 llodvth = 0
+ wlodvth = 1 lku0 = 0 wku0 = 0
+ pku0 = 0 lkvth0 = 0 wkvth0 = 7.3E-7
+ pkvth0 = 0 stk2 = 0 lodk2 = 1
+ steta0 = 0 lodeta0 = 1

.model plowvt_model.18 pmos
+ level = 54 lmin = 1.5E-6 lmax = 2E-6 wmin = 3E-6
+ wmax = 5E-6 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 4.23E-9
+ toxm = 4.23E-9 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 9.999999999999999E22 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {7.476E-9+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {2.8E-9-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = -7.916E-9 dwb = 0 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = -0.438272581967641 lvth0 = -3.365680408303202E-8
+ wvth0 = 1.583097125442938E-7 pvth0 = -4.625770650022766E-14 k1 = 0.64774
+ k2 = -0.05250534235076 lk2 = 9.840997767313542E-9 wk2 = 4.821266018031074E-8
+ pk2 = -9.174371204829791E-14 k3 = 3.39 k3b = 1
+ w0 = 1E-8 lpe0 = 0 lpeb = 0
+ vbm = -3 dvtp0 = 0 dvtp1 = 0
+ dvt0 = 2.4422 dvt1 = 0.16136 dvt2 = 0.026237
+ dvt0w = 0.5 dvt1w = 1.9281E6 dvt2w = -0.032
+ vfbsdoff = 0 u0 = 1.919212886664862E-3 lu0 = 1.02003340750869E-9
+ wu0 = 1.78546059096779E-9 pu0 = -2.540404054010693E-15 ua = -3.003633671472641E-9
+ lua = -4.130410962504846E-16 wua = 3.43082526162064E-16 pua = 1.232947498280317E-21
+ ub = 2.892636887468803E-18 lub = 9.434571802843813E-25 wub = 8.84503313502497E-27
+ pub = -2.816264969093532E-30 uc = -3.342407413682558E-11 luc = 1.92970422953285E-16
+ wuc = 2.52550207341983E-16 puc = -5.760259750958574E-22 ud = 0
+ up = 0 lp = 1 eu = 1.67
+ vsat = 5.199177924737537E5 lvsat = -0.790097101309654 wvsat = -1.182550026108194
+ pvsat = 2.358477772070182E-6 a0 = 1.83259450571751 la0 = 4.009081076545377E-7
+ wa0 = 9.818426055422684E-8 pa0 = -2.952997959640246E-12 ags = -0.130137004887424
+ lags = 1.526883444072982E-6 wags = 1.074878187784394E-6 pags = -3.476867594521075E-12
+ b0 = 0 b1 = 2.1073E-24 keta = -0.01258
+ a1 = 0 a2 = 0.46703705 rdsw = 484.7
+ rdswmin = 0 rdw = 0 rdwmin = 0
+ rsw = 0 rswmin = 0 prwb = 0.1
+ prwg = 0.052 wr = 1 voff = -0.1819
+ voffl = 0 minv = 0 nfactor = 2.5373
+ eta0 = 0.2 etab = -2.5E-4 dsub = 1
+ cit = -6.393105E-11 cdsc = 2.8125E-7 cdscb = 1E-4
+ cdscd = 1E-10 pclm = 0.030097 pdiblc1 = 0
+ pdiblc2 = -7.423973214826881E-3 lpdiblc2 = 2.967777192122674E-8 wpdiblc2 = 2.761692790802024E-8
+ ppdiblc2 = -6.097768040955457E-14 pdiblcb = -0.025 drout = 0.43496
+ pscbe1 = 8E8 pscbe2 = 8.6797E-9 pvag = 0
+ delta = -0.014403468893824 ldelta = 6.22313738928379E-8 wdelta = 2.031245788404278E-7
+ pdelta = -2.669907891959552E-13 fprout = 0 pdits = 0
+ pditsl = 0 pditsd = 0 lambda = 0
+ vtl = 0 lc = 5E-9 xn = 3
+ alpha0 = 5.0449517E-13 alpha1 = -4.0583656E-18 beta0 = 6.2016506
+ aigbacc = 0.43 bigbacc = 0.054 cigbacc = 0.075
+ nigbacc = 1 aigbinv = 0.35 bigbinv = 0.03
+ cigbinv = 6E-3 eigbinv = 1.1 nigbinv = 3
+ aigc = 0.43 bigc = 0.054 cigc = 0.075
+ aigsd = 0.43 bigsd = 0.054 cigsd = 0.075
+ dlcig = 0 nigc = 1 poxedge = 1
+ pigcd = 1 ntox = 1 toxref = 4.23E-9
+ agidl = 0 bgidl = 2.3E9 cgidl = 0.5
+ egidl = 0.8 noia = 3E41 noib = 0
+ noic = 0 em = 4.1E7 af = 1
+ ef = 0.88 kf = 0 lintnoi = 0
+ tnoia = 2.5E7 tnoib = 0 ntnoi = 1
+ rnoia = 0.69 rnoib = 0.34 xpart = 0
+ cgso = {2E-11/sw_func_tox_lv_ratio} cgdo = {2E-11/sw_func_tox_lv_ratio} cgbo = {1E-13/sw_func_tox_lv_ratio}
+ ckappas = 0.6 cf = 0 clc = 7E-8
+ cle = 0.492 dlc = -1.2E-8 dwc = 0
+ vfbcv = -1 noff = 2.6123 voffcv = 0.112
+ acde = 0.44 moin = 8.7 cgsl = {0/sw_func_tox_lv_ratio}
+ cgdl = {0/sw_func_tox_lv_ratio} ijthsrev = 0.1 ijthsfwd = 0.1
+ xjbvs = 1 bvs = 12.69 jss = 2.1483E-5
+ jsws = 1.4472E-10 cjs = {7.682E-04*sw_func_psd_nw_cj} mjs = 0.3362
+ mjsws = 0.2659 cjsws = {9.160236799999998E-11*sw_func_psd_nw_cj} cjswgs = {2.39155046E-10*sw_func_psd_nw_cj}
+ mjswgs = 0.9274 pbs = 0.6587 pbsws = 0.7418
+ pbswgs = 1.4338 xrcrg1 = 12 xrcrg2 = 1
+ rbpb = 50 rbpd = 50 rbps = 50
+ rbdb = 50 rbsb = 50 gbmin = 1E-12
+ tnom = 30 ute = -0.13298 kt1 = -0.367860328064001
+ lkt1 = -4.457278017091573E-7 wkt1 = -6.671273982332113E-7 pkt1 = 1.330518883036317E-12
+ kt1l = 0 kt2 = 0.096682138277351 lkt2 = -3.026046045803479E-7
+ wkt2 = -4.529127906605287E-7 pkt2 = 9.032892696933584E-13 ua1 = 9.090011607976962E-10
+ lua1 = -4.246300190949253E-16 wua1 = -6.355500347168415E-16 pua1 = 1.267540989239269E-21
+ ub1 = -9.483448068193279E-19 lub1 = 1.648301410720468E-24 wub1 = 2.467037118666422E-24
+ pub1 = -4.920258829468312E-30 uc1 = -9.961E-12 at = 1.110114556206656E6
+ lat = -1.698221833197147 wat = -2.404237026273103 pat = 4.684756987170884E-6
+ prt = 0 njs = 1.3632 xtis = 5.2
+ tpb = 1.671E-3 tpbsw = 1.246E-3 tpbswg = 0
+ tcj = 1.2407E-3 tcjsw = 3.7357E-4 tcjswg = 2E-12
+ tvoff = 0 tvfbsdoff = 0 saref = 3E-6
+ sbref = 3E-6 wlod = 0 ku0 = 5.9E-8
+ kvsat = 0 kvth0 = 1.76E-8 tku0 = 0
+ llodku0 = 0 wlodku0 = 1 llodvth = 0
+ wlodvth = 1 lku0 = 0 wku0 = 0
+ pku0 = 0 lkvth0 = 0 wkvth0 = 7.3E-7
+ pkvth0 = 0 stk2 = 0 lodk2 = 1
+ steta0 = 0 lodeta0 = 1

.model plowvt_model.19 pmos
+ level = 54 lmin = 1E-6 lmax = 1.5E-6 wmin = 3E-6
+ wmax = 5E-6 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 4.23E-9
+ toxm = 4.23E-9 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 9.999999999999999E22 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {7.476E-9+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {2.8E-9-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = -7.916E-9 dwb = 0 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = -0.483828760510342 lvth0 = 3.442234913118033E-8
+ wvth0 = 2.738783083578538E-7 pvth0 = -2.189634160840115E-13 k1 = 0.64774
+ k2 = -0.038865798427978 lk2 = -1.054193667089247E-8 wk2 = -5.26460091158637E-8
+ pk2 = 5.897948334790517E-14 k3 = 3.39 k3b = 1
+ w0 = 1E-8 lpe0 = 0 lpeb = 0
+ vbm = -3 dvtp0 = 0 dvtp1 = 0
+ dvt0 = 2.4422 dvt1 = 0.16136 dvt2 = 0.026237
+ dvt0w = 0.5 dvt1w = 1.9281E6 dvt2w = -0.032
+ vfbsdoff = 0 u0 = 3.556774614033156E-3 lu0 = -1.427138837870488E-9
+ wu0 = -7.087228491307668E-9 pu0 = 1.071894251054175E-14 ua = -3.161590541528959E-9
+ lua = -1.769903496383235E-16 wua = 1.811493737718542E-16 pua = 1.474940401212246E-21
+ ub = 3.631122075896321E-18 lub = -1.601350853017013E-25 wub = -2.409882252602801E-24
+ pub = 7.982810867130755E-31 uc = 1.588360267414017E-10 luc = -9.434307179913781E-17
+ wuc = -5.153121542444381E-16 puc = 5.714675380588901E-22 ud = 0
+ up = 0 lp = 1 eu = 1.67
+ vsat = -2.950518844853378E5 lvsat = 0.427793583938012 wvsat = 1.250173578159189
+ pvsat = -1.276984382146995E-6 a0 = 2.670256878585164 la0 = -8.508945423588857E-7
+ wa0 = -2.676230509259168E-6 pa0 = 1.193087472368891E-12 ags = 1.218875402735277
+ lags = -4.890806978783813E-7 wags = -2.608836892356228E-6 pags = 2.028076221241071E-12
+ b0 = 0 b1 = 2.1073E-24 keta = -0.01258
+ a1 = 0 a2 = 0.46703705 rdsw = 484.7
+ rdswmin = 0 rdw = 0 rdwmin = 0
+ rsw = 0 rswmin = 0 prwb = 0.1
+ prwg = 0.052 wr = 1 voff = -0.1819
+ voffl = 0 minv = 0 nfactor = 6.773703046768642
+ lnfactor = -6.330880713091057E-6 wnfactor = -2.111867253548793E-5 pnfactor = 3.155974423703315E-11
+ eta0 = 0.2 etab = -2.5E-4 dsub = 1
+ cit = -6.393105E-11 cdsc = 2.8125E-7 cdscb = 1E-4
+ cdscd = 1E-10 pclm = 0.030097 pdiblc1 = 0
+ pdiblc2 = -0.014835746674623 lpdiblc2 = 4.075392617954564E-8 wpdiblc2 = 4.334727887501064E-8
+ ppdiblc2 = -8.448511689462502E-14 pdiblcb = -0.025 drout = 0.43496
+ pscbe1 = 8E8 pscbe2 = 8.6797E-9 pvag = 0
+ delta = 0.037745694016467 ldelta = -1.570033516030138E-8 wdelta = -1.276670773680706E-7
+ pdelta = 2.273442618420248E-13 fprout = 0 pdits = 0
+ pditsl = 0 pditsd = 0 lambda = 0
+ vtl = 0 lc = 5E-9 xn = 3
+ alpha0 = 5.0449517E-13 alpha1 = -4.0583656E-18 beta0 = 6.2016506
+ aigbacc = 0.43 bigbacc = 0.054 cigbacc = 0.075
+ nigbacc = 1 aigbinv = 0.35 bigbinv = 0.03
+ cigbinv = 6E-3 eigbinv = 1.1 nigbinv = 3
+ aigc = 0.43 bigc = 0.054 cigc = 0.075
+ aigsd = 0.43 bigsd = 0.054 cigsd = 0.075
+ dlcig = 0 nigc = 1 poxedge = 1
+ pigcd = 1 ntox = 1 toxref = 4.23E-9
+ agidl = 0 bgidl = 2.3E9 cgidl = 0.5
+ egidl = 0.8 noia = 3E41 noib = 0
+ noic = 0 em = 4.1E7 af = 1
+ ef = 0.88 kf = 0 lintnoi = 0
+ tnoia = 2.5E7 tnoib = 0 ntnoi = 1
+ rnoia = 0.69 rnoib = 0.34 xpart = 0
+ cgso = {2E-11/sw_func_tox_lv_ratio} cgdo = {2E-11/sw_func_tox_lv_ratio} cgbo = {1E-13/sw_func_tox_lv_ratio}
+ ckappas = 0.6 cf = 0 clc = 7E-8
+ cle = 0.492 dlc = -1.2E-8 dwc = 0
+ vfbcv = -1 noff = 2.6123 voffcv = 0.112
+ acde = 0.44 moin = 8.7 cgsl = {0/sw_func_tox_lv_ratio}
+ cgdl = {0/sw_func_tox_lv_ratio} ijthsrev = 0.1 ijthsfwd = 0.1
+ xjbvs = 1 bvs = 12.69 jss = 2.1483E-5
+ jsws = 1.4472E-10 cjs = {7.682E-04*sw_func_psd_nw_cj} mjs = 0.3362
+ mjsws = 0.2659 cjsws = {9.160236799999998E-11*sw_func_psd_nw_cj} cjswgs = {2.39155046E-10*sw_func_psd_nw_cj}
+ mjswgs = 0.9274 pbs = 0.6587 pbsws = 0.7418
+ pbswgs = 1.4338 xrcrg1 = 12 xrcrg2 = 1
+ rbpb = 50 rbpd = 50 rbps = 50
+ rbdb = 50 rbsb = 50 gbmin = 1E-12
+ tnom = 30 ute = -0.669196296617409 lute = 8.013216336650553E-7
+ wute = 3.042172005725171E-6 pute = -4.546221845355695E-12 kt1 = -0.854318306559999
+ lkt1 = 2.81235001355263E-7 wkt1 = 9.630729214323121E-7 pkt1 = -1.105652474671841E-12
+ kt1l = 0 kt2 = -0.245088359077351 lkt2 = 2.081372266665174E-7
+ wkt2 = 4.529127906605287E-7 pkt2 = -4.503764790328297E-13 ua1 = 5.918468712023039E-10
+ lua1 = 4.932535127642901E-17 wua1 = 6.355500347168416E-16 pua1 = -6.319909545224272E-22
+ ub1 = 4.839473348193283E-19 lub1 = -4.921159657443398E-25 wub1 = -2.467037118666422E-24
+ pub1 = 2.45322171080189E-30 uc1 = -9.961E-12 at = -6.458038850709765E5
+ lat = 0.925822685448147 wat = 2.772365995859732 pat = -3.051158569104424E-6
+ prt = 0 njs = 1.3632 xtis = 5.2
+ tpb = 1.671E-3 tpbsw = 1.246E-3 tpbswg = 0
+ tcj = 1.2407E-3 tcjsw = 3.7357E-4 tcjswg = 2E-12
+ tvoff = 0 tvfbsdoff = 0 saref = 3E-6
+ sbref = 3E-6 wlod = 0 ku0 = 5.9E-8
+ kvsat = 0 kvth0 = 1.76E-8 tku0 = 0
+ llodku0 = 0 wlodku0 = 1 llodvth = 0
+ wlodvth = 1 lku0 = 0 wku0 = 0
+ pku0 = 0 lkvth0 = 0 wkvth0 = 7.3E-7
+ pkvth0 = 0 stk2 = 0 lodk2 = 1
+ steta0 = 0 lodeta0 = 1

.model plowvt_model.20 pmos
+ level = 54 lmin = 5E-7 lmax = 1E-6 wmin = 3E-6
+ wmax = 5E-6 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 4.23E-9
+ toxm = 4.23E-9 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 9.999999999999999E22 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {7.476E-9+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {2.8E-9-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = -7.916E-9 dwb = 0 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = -0.421165091610874 lvth0 = -2.789040322245127E-8
+ wvth0 = -6.474339260058142E-8 pvth0 = 1.177620033490564E-13 k1 = 0.64774
+ k2 = -0.042174041795666 lk2 = -7.252219466063404E-9 wk2 = -1.047399276916289E-8
+ pk2 = 1.704363029274588E-14 k3 = 3.39 k3b = 1
+ w0 = 1E-8 lpe0 = 0 lpeb = 0
+ vbm = -3 dvtp0 = 0 dvtp1 = 0
+ dvt0 = 2.4422 dvt1 = 0.16136 dvt2 = 0.026237
+ dvt0w = 0.5 dvt1w = 1.9281E6 dvt2w = -0.032
+ vfbsdoff = 0 u0 = 7.659748549211749E-4 lu0 = 1.348032442590465E-9
+ wu0 = 8.395580388005153E-9 pu0 = -4.677162639046919E-15 ua = -3.860260525176961E-9
+ lua = 5.17767082101249E-16 wua = 3.307207888030434E-15 pua = -1.633612185366485E-21
+ ub = 4.002440453939199E-18 lub = -5.293740804275401E-25 wub = -3.1962116505503E-24
+ pub = 1.580207040032068E-30 uc = 7.475688873712637E-11 luc = -1.073477696768647E-17
+ wuc = 8.348977963130966E-17 puc = -2.398110498715342E-23 ud = 0
+ up = 0 lp = 1 eu = 1.67
+ vsat = 1.809084120261633E4 lvsat = 0.11640445751391 wvsat = 0.334224579040561
+ pvsat = -3.66164697423431E-7 a0 = 1.71406973730811 la0 = 9.993795092701787E-8
+ wa0 = -1.918386879800898E-6 pa0 = 4.394877672355871E-13 ags = 1.057449275384275
+ lags = -3.285585568405457E-7 wags = -8.755440330156967E-7 pags = 3.044898019128462E-13
+ b0 = 1.43666401937664E-6 lb0 = -1.428618700868131E-12 wb0 = -1.046161472265801E-12
+ pb0 = 1.040302968021113E-18 b1 = 2.1073E-24 keta = -0.01258
+ a1 = 0 a2 = 0.46703705 rdsw = 484.7
+ rdswmin = 0 rdw = 0 rdwmin = 0
+ rsw = 0 rswmin = 0 prwb = 0.1
+ prwg = 0.052 wr = 1 voff = -0.1819
+ voffl = 0 minv = 0 nfactor = 0.407169747199999
+ wnfactor = 1.061880155646014E-5 eta0 = 0.2 etab = -2.5E-4
+ dsub = 1 cit = -6.393105E-11 cdsc = 2.8125E-7
+ cdscb = 1E-4 cdscd = 1E-10 pclm = 0.030097
+ pdiblc1 = 0 pdiblc2 = -9.80418428401279E-3 lpdiblc2 = 3.575054053832312E-8
+ wpdiblc2 = -2.694381612464978E-8 ppdiblc2 = -1.45876520269627E-14 pdiblcb = -0.025
+ drout = 0.43496 pscbe1 = 8E8 pscbe2 = 8.6797E-9
+ pvag = 0 delta = 2.953963186822409E-3 ldelta = 1.889656197669739E-8
+ wdelta = 1.263243227685646E-7 pdelta = -2.52247864538452E-14 fprout = 0
+ pdits = 0 pditsl = 0 pditsd = 0
+ lambda = 0 vtl = 0 lc = 5E-9
+ xn = 3 alpha0 = 5.0449517E-13 alpha1 = -4.0583656E-18
+ beta0 = 6.2016506 aigbacc = 0.43 bigbacc = 0.054
+ cigbacc = 0.075 nigbacc = 1 aigbinv = 0.35
+ bigbinv = 0.03 cigbinv = 6E-3 eigbinv = 1.1
+ nigbinv = 3 aigc = 0.43 bigc = 0.054
+ cigc = 0.075 aigsd = 0.43 bigsd = 0.054
+ cigsd = 0.075 dlcig = 0 nigc = 1
+ poxedge = 1 pigcd = 1 ntox = 1
+ toxref = 4.23E-9 agidl = 0 bgidl = 2.3E9
+ cgidl = 0.5 egidl = 0.8 noia = 3E41
+ noib = 0 noic = 0 em = 4.1E7
+ af = 1 ef = 0.88 kf = 0
+ lintnoi = 0 tnoia = 2.5E7 tnoib = 0
+ ntnoi = 1 rnoia = 0.69 rnoib = 0.34
+ xpart = 0 cgso = {2E-11/sw_func_tox_lv_ratio} cgdo = {2E-11/sw_func_tox_lv_ratio}
+ cgbo = {1E-13/sw_func_tox_lv_ratio} ckappas = 0.6 cf = 0
+ clc = 7E-8 cle = 0.492 dlc = -1.2E-8
+ dwc = 0 vfbcv = -1 noff = 2.6123
+ voffcv = 0.112 acde = 0.44 moin = 8.7
+ cgsl = {0/sw_func_tox_lv_ratio} cgdl = {0/sw_func_tox_lv_ratio} ijthsrev = 0.1
+ ijthsfwd = 0.1 xjbvs = 1 bvs = 12.69
+ jss = 2.1483E-5 jsws = 1.4472E-10 cjs = {7.682E-04*sw_func_psd_nw_cj}
+ mjs = 0.3362 mjsws = 0.2659 cjsws = {9.160236799999998E-11*sw_func_psd_nw_cj}
+ cjswgs = {2.39155046E-10*sw_func_psd_nw_cj} mjswgs = 0.9274 pbs = 0.6587
+ pbsws = 0.7418 pbswgs = 1.4338 xrcrg1 = 12
+ xrcrg2 = 1 rbpb = 50 rbpd = 50
+ rbps = 50 rbdb = 50 rbsb = 50
+ gbmin = 1E-12 tnom = 30 ute = 0.612840231376576
+ lute = -4.735354897721632E-7 wute = -2.778350976221291E-6 pute = 1.241706207891866E-12
+ kt1 = -0.534983136 lkt1 = -3.631189224959974E-8 wkt1 = -1.488060756230385E-7
+ kt1l = 0 kt2 = -8.330096427020789E-3 lkt2 = -2.729518971297053E-8
+ wkt2 = -3.708649776154645E-8 pkt2 = 3.687881337408179E-14 ua1 = 3.8940488E-10
+ lua1 = 2.50633667328E-16 ub1 = 5.1769597606336E-19 lub1 = -5.256756145974052E-25
+ wub1 = 2.644831570179714E-25 pub1 = -2.630020513386707E-31 uc1 = -2.284941472E-11
+ luc1 = 1.2816239597568E-17 at = 5.13853042990208E5 lat = -0.227340163815895
+ wat = -0.614826467311553 pat = 3.170656162731013E-7 prt = 0
+ njs = 1.3632 xtis = 5.2 tpb = 1.671E-3
+ tpbsw = 1.246E-3 tpbswg = 0 tcj = 1.2407E-3
+ tcjsw = 3.7357E-4 tcjswg = 2E-12 tvoff = 0
+ tvfbsdoff = 0 saref = 2.74E-6 sbref = 2.74E-6
+ wlod = 0 ku0 = 5.9E-8 kvsat = 0
+ kvth0 = 1.76E-8 tku0 = 0 llodku0 = 0
+ wlodku0 = 1 llodvth = 0 wlodvth = 1
+ lku0 = 0 wku0 = 0 pku0 = 0
+ lkvth0 = 0 wkvth0 = 7.3E-7 pkvth0 = 0
+ stk2 = 0 lodk2 = 1 steta0 = 0
+ lodeta0 = 1

.model plowvt_model.21 pmos
+ level = 54 lmin = 3.5E-7 lmax = 5E-7 wmin = 3E-6
+ wmax = 5E-6 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 4.23E-9
+ toxm = 4.23E-9 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 9.999999999999999E22 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {7.476E-9+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {2.8E-9-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = -7.916E-9 dwb = 0 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = -0.407798362851808 lvth0 = -3.449891392093337E-8
+ wvth0 = -1.848320860538086E-7 pvth0 = 1.771338533923319E-13 k1 = 0.64774
+ k2 = -0.050056874402566 lk2 = -3.354947025212181E-9 wk2 = -9.307529679806387E-8
+ pk2 = 5.788171500463453E-14 k3 = 3.39 k3b = 1
+ w0 = 1E-8 lpe0 = 0 lpeb = 0
+ vbm = -3 dvtp0 = 0 dvtp1 = 0
+ dvt0 = 2.4422 dvt1 = 0.16136 dvt2 = 0.026237
+ dvt0w = 0.5 dvt1w = 1.9281E6 dvt2w = -0.032
+ vfbsdoff = 0 u0 = 2.516996828581534E-3 lu0 = 4.823271788127838E-10
+ wu0 = 1.55267931839027E-9 pu0 = -1.294032350229321E-15 ua = -2.883571214224001E-9
+ lua = 3.489188676610616E-17 wua = 1.17315733899693E-15 pua = -5.785375939243209E-22
+ ub = 2.725739066796801E-18 lub = 1.018270853756615E-25 wub = -1.609212710759659E-24
+ pub = 7.955947641995753E-31 uc = -1.338483518969599E-11 luc = 3.284249134173449E-17
+ wuc = 3.309291173089157E-16 puc = -1.463151135349618E-22 ud = 0
+ up = 0 lp = 1 eu = 1.67
+ vsat = 6.576482278432767E5 lvsat = -0.199792714441232 wvsat = -1.650280235319073
+ pvsat = 6.149744827959719E-7 a0 = 5.712683401723647 la0 = -1.876976644760024E-6
+ wa0 = -1.183205582345986E-5 pa0 = 5.340805692980576E-12 ags = -0.11421133096544
+ lags = 2.507104469387536E-7 wags = 1.254052488275726E-6 pags = -7.483827182136328E-13
+ b0 = -4.788880064588801E-6 lb0 = 1.649290294244383E-12 wb0 = 3.487204907552672E-12
+ pb0 = -1.20099337016114E-18 b1 = 2.1073E-24 keta = -0.01258
+ a1 = 0 a2 = 0.46703705 rdsw = 484.7
+ rdswmin = 0 rdw = 0 rdwmin = 0
+ rsw = 0 rswmin = 0 prwb = 0.1
+ prwg = 0.052 wr = 1 voff = -0.1819
+ voffl = 0 minv = 0 nfactor = 0.407169747199999
+ wnfactor = 1.061880155646014E-5 eta0 = 0.2 etab = -2.5E-4
+ dsub = 1 cit = -6.393105E-11 cdsc = 2.8125E-7
+ cdscb = 1E-4 cdscd = 1E-10 pclm = 0.030097
+ pdiblc1 = 0 pdiblc2 = -0.030977732212064 lpdiblc2 = 4.621874263395164E-8
+ wpdiblc2 = -1.484241201881308E-7 ppdiblc2 = 4.547221030202232E-14 pdiblcb = -0.025
+ drout = 0.43496 pscbe1 = 8E8 pscbe2 = 8.6797E-9
+ pvag = 0 delta = 0.059235897445824 ldelta = -8.929226320952972E-9
+ wdelta = -1.24242478152654E-7 pdelta = 9.865543992160523E-14 fprout = 0
+ pdits = 0 pditsl = 0 pditsd = 0
+ lambda = 0 vtl = 0 lc = 5E-9
+ xn = 3 alpha0 = 5.0449517E-13 alpha1 = -4.0583656E-18
+ beta0 = 6.2016506 aigbacc = 0.43 bigbacc = 0.054
+ cigbacc = 0.075 nigbacc = 1 aigbinv = 0.35
+ bigbinv = 0.03 cigbinv = 6E-3 eigbinv = 1.1
+ nigbinv = 3 aigc = 0.43 bigc = 0.054
+ cigc = 0.075 aigsd = 0.43 bigsd = 0.054
+ cigsd = 0.075 dlcig = 0 nigc = 1
+ poxedge = 1 pigcd = 1 ntox = 1
+ toxref = 4.23E-9 agidl = 0 bgidl = 2.3E9
+ cgidl = 0.5 egidl = 0.8 noia = 3E41
+ noib = 0 noic = 0 em = 4.1E7
+ af = 1 ef = 0.88 kf = 0
+ lintnoi = 0 tnoia = 2.5E7 tnoib = 0
+ ntnoi = 1 rnoia = 0.69 rnoib = 0.34
+ xpart = 0 cgso = {2E-11/sw_func_tox_lv_ratio} cgdo = {2E-11/sw_func_tox_lv_ratio}
+ cgbo = {1E-13/sw_func_tox_lv_ratio} ckappas = 0.6 cf = 0
+ clc = 7E-8 cle = 0.492 dlc = -1.2E-8
+ dwc = 0 vfbcv = -1 noff = 2.6123
+ voffcv = 0.112 acde = 0.44 moin = 8.7
+ cgsl = {0/sw_func_tox_lv_ratio} cgdl = {0/sw_func_tox_lv_ratio} ijthsrev = 0.1
+ ijthsfwd = 0.1 xjbvs = 1 bvs = 12.69
+ jss = 2.1483E-5 jsws = 1.4472E-10 cjs = {7.682E-04*sw_func_psd_nw_cj}
+ mjs = 0.3362 mjsws = 0.2659 cjsws = {9.160236799999998E-11*sw_func_psd_nw_cj}
+ cjswgs = {2.39155046E-10*sw_func_psd_nw_cj} mjswgs = 0.9274 pbs = 0.6587
+ pbsws = 0.7418 pbswgs = 1.4338 xrcrg1 = 12
+ xrcrg2 = 1 rbpb = 50 rbpd = 50
+ rbps = 50 rbdb = 50 rbsb = 50
+ gbmin = 1E-12 tnom = 30 ute = -0.22207178253056
+ lute = -6.075499009647515E-8 wute = -8.794034316795974E-7 pute = 3.028665418704533E-13
+ kt1 = -0.68016859104 lkt1 = 3.546779672217601E-8 wkt1 = 2.202329919220994E-8
+ pkt1 = -8.445804290865966E-14 kt1l = 0 kt2 = -0.080813489243264
+ lkt2 = 8.54059969538013E-9 wkt2 = 1.236216592051548E-7 pkt2 = -4.257529943025533E-14
+ ua1 = 8.9635E-10 ub1 = -4.223690402112E-19 lub1 = -6.090747055126271E-26
+ wub1 = -8.816105233932379E-25 pub1 = 3.036266642566311E-31 uc1 = 3.0734E-12
+ at = 1.2016489758976E5 lat = -0.032700744729913 wat = 0.08730273889513
+ pat = -3.006706327548281E-8 prt = 0 njs = 1.3632
+ xtis = 5.2 tpb = 1.671E-3 tpbsw = 1.246E-3
+ tpbswg = 0 tcj = 1.2407E-3 tcjsw = 3.7357E-4
+ tcjswg = 2E-12 tvoff = 0 tvfbsdoff = 0
+ saref = 1.74E-6 sbref = 1.74E-6 wlod = 0
+ ku0 = 5.9E-8 kvsat = 0 kvth0 = 1.76E-8
+ tku0 = 0 llodku0 = 0 wlodku0 = 1
+ llodvth = 0 wlodvth = 1 lku0 = 0
+ wku0 = 0 pku0 = 0 lkvth0 = 0
+ wkvth0 = 7.3E-7 pkvth0 = 0 stk2 = 0
+ lodk2 = 1 steta0 = 0 lodeta0 = 1

.model plowvt_model.22 pmos
+ level = 54 lmin = 8E-6 lmax = 2.02E-5 wmin = 1E-6
+ wmax = 3E-6 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 4.23E-9
+ toxm = 4.23E-9 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 9.999999999999999E22 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {7.476E-9+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {2.8E-9-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = -7.916E-9 dwb = 0 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = -0.4499316647968 wvth0 = 4.525770016875826E-8
+ k1 = 0.64774 k2 = -0.0509446978492 wk2 = 1.210466172455876E-8
+ k3 = 3.39 k3b = 1 w0 = 1E-8
+ lpe0 = 0 lpeb = 0 vbm = -3
+ dvtp0 = 0 dvtp1 = 0 dvt0 = 2.4422
+ dvt1 = 0.16136 dvt2 = 0.026237 dvt0w = 0.5
+ dvt1w = 1.9281E6 dvt2w = -0.032 vfbsdoff = 0
+ u0 = 2.832952674432E-3 wu0 = -2.716473513078928E-10 ua = -2.8451063376E-9
+ wua = -4.057773475979487E-17 ub = 2.8737319344E-18 wub = 6.527722548314926E-26
+ uc = 5.9129332256E-11 wuc = 5.375079647891704E-18 ud = 0
+ up = 0 lp = 1 eu = 1.67
+ vsat = 1.2376E5 a0 = 1.87941253692 wa0 = -3.989114772599722E-7
+ ags = 0.39855725812 wags = -1.214832689565898E-7 b0 = 0
+ b1 = 2.1073E-24 keta = -0.01258 a1 = 0
+ a2 = 0.46703705 rdsw = 484.7 rdswmin = 0
+ rdw = 0 rdwmin = 0 rsw = 0
+ rswmin = 0 prwb = 0.1 prwg = 0.052
+ wr = 1 voff = -0.1819 voffl = 0
+ minv = 0 nfactor = 2.5373 eta0 = 0.2
+ etab = -2.5E-4 dsub = 1 cit = -6.393105E-11
+ cdsc = 2.8125E-7 cdscb = 1E-4 cdscd = 1E-10
+ pclm = 0.030097 pdiblc1 = 0 pdiblc2 = 2.6689050296E-3
+ wpdiblc2 = -1.257615735997421E-9 pdiblcb = -0.025 drout = 0.43496
+ pscbe1 = 8E8 pscbe2 = 8.6797E-9 pvag = 0
+ delta = 0.02448898624 wdelta = -1.140881238173952E-8 fprout = 0
+ pdits = 0 pditsl = 0 pditsd = 0
+ lambda = 0 vtl = 0 lc = 5E-9
+ xn = 3 alpha0 = 5.0449517E-13 alpha1 = -4.0583656E-18
+ beta0 = 6.2016506 aigbacc = 0.43 bigbacc = 0.054
+ cigbacc = 0.075 nigbacc = 1 aigbinv = 0.35
+ bigbinv = 0.03 cigbinv = 6E-3 eigbinv = 1.1
+ nigbinv = 3 aigc = 0.43 bigc = 0.054
+ cigc = 0.075 aigsd = 0.43 bigsd = 0.054
+ cigsd = 0.075 dlcig = 0 nigc = 1
+ poxedge = 1 pigcd = 1 ntox = 1
+ toxref = 4.23E-9 agidl = 0 bgidl = 2.3E9
+ cgidl = 0.5 egidl = 0.8 noia = 3E41
+ noib = 0 noic = 0 em = 4.1E7
+ af = 1 ef = 0.88 kf = 0
+ lintnoi = 0 tnoia = 2.5E7 tnoib = 0
+ ntnoi = 1 rnoia = 0.69 rnoib = 0.34
+ xpart = 0 cgso = {2E-11/sw_func_tox_lv_ratio} cgdo = {2E-11/sw_func_tox_lv_ratio}
+ cgbo = {1E-13/sw_func_tox_lv_ratio} ckappas = 0.6 cf = 0
+ clc = 7E-8 cle = 0.492 dlc = -1.2E-8
+ dwc = 0 vfbcv = -1 noff = 2.6123
+ voffcv = 0.112 acde = 0.44 moin = 8.7
+ cgsl = {0/sw_func_tox_lv_ratio} cgdl = {0/sw_func_tox_lv_ratio} ijthsrev = 0.1
+ ijthsfwd = 0.1 xjbvs = 1 bvs = 12.69
+ jss = 2.1483E-5 jsws = 1.4472E-10 cjs = {7.682E-04*sw_func_psd_nw_cj}
+ mjs = 0.3362 mjsws = 0.2659 cjsws = {9.160236799999998E-11*sw_func_psd_nw_cj}
+ cjswgs = {2.39155046E-10*sw_func_psd_nw_cj} mjswgs = 0.9274 pbs = 0.6587
+ pbsws = 0.7418 pbswgs = 1.4338 xrcrg1 = 12
+ xrcrg2 = 1 rbpb = 50 rbpd = 50
+ rbps = 50 rbdb = 50 rbsb = 50
+ gbmin = 1E-12 tnom = 30 ute = -0.29175
+ kt1 = -0.59149952 wkt1 = -2.940415562303986E-8 kt1l = 0
+ kt2 = -0.055045 ua1 = 6.8217E-10 ub1 = -1.5013E-19
+ uc1 = -9.961E-12 at = 2.8691660352E5 wat = -0.012467361984169
+ prt = 0 njs = 1.3632 xtis = 5.2
+ tpb = 1.671E-3 tpbsw = 1.246E-3 tpbswg = 0
+ tcj = 1.2407E-3 tcjsw = 3.7357E-4 tcjswg = 2E-12
+ tvoff = 0 tvfbsdoff = 0 saref = 3E-6
+ sbref = 3E-6 wlod = 0 ku0 = 5.9E-8
+ kvsat = 0 kvth0 = 1.76E-8 tku0 = 0
+ llodku0 = 0 wlodku0 = 1 llodvth = 0
+ wlodvth = 1 lku0 = 0 wku0 = 0
+ pku0 = 0 lkvth0 = 0 wkvth0 = 7.3E-7
+ pkvth0 = 0 stk2 = 0 lodk2 = 1
+ steta0 = 0 lodeta0 = 1

.model plowvt_model.23 pmos
+ level = 54 lmin = 4E-6 lmax = 8E-6 wmin = 1E-6
+ wmax = 3E-6 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 4.23E-9
+ toxm = 4.23E-9 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 9.999999999999999E22 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {7.476E-9+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {2.8E-9-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = -7.916E-9 dwb = 0 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = -0.470384023483016 lvth0 = 1.635043362810881E-7
+ wvth0 = 5.126066980452684E-8 pvth0 = -4.799014045618833E-14 k1 = 0.64774
+ k2 = -0.056175001290615 lk2 = 4.181313783204959E-8 wk2 = 1.569135092925999E-8
+ pk2 = -2.867342817806351E-14 k3 = 3.39 k3b = 1
+ w0 = 1E-8 lpe0 = 0 lpeb = 0
+ vbm = -3 dvtp0 = 0 dvtp1 = 0
+ dvt0 = 2.4422 dvt1 = 0.16136 dvt2 = 0.026237
+ dvt0w = 0.5 dvt1w = 1.9281E6 dvt2w = -0.032
+ vfbsdoff = 0 u0 = 3.037702043719614E-3 lu0 = -1.636848357832901E-9
+ wu0 = -4.804167406731458E-10 pu0 = 1.668986006341578E-15 ua = -2.824985026928E-9
+ lua = -1.608578060362379E-16 wua = -1.121474495462723E-17 pua = -2.347394856984321E-22
+ ub = 2.9145541951112E-18 lub = -3.263494810296166E-25 wub = -5.657918220829666E-26
+ pub = 9.741688656484952E-31 uc = 5.9129332256E-11 wuc = 5.375079647891704E-18
+ ud = 0 up = 0 lp = 1
+ eu = 1.67 vsat = 1.2376E5 a0 = 1.858357855766645
+ la0 = 1.683195430123828E-7 wa0 = -4.702371157957053E-7 pa0 = 5.70205684710065E-13
+ ags = 0.365866956477119 lags = 2.613393474538461E-7 wags = -1.377107252724158E-7
+ pags = 1.297287767712394E-13 b0 = 0 b1 = 2.1073E-24
+ keta = -0.01258 a1 = 0 a2 = 0.46703705
+ rdsw = 484.7 rdswmin = 0 rdw = 0
+ rdwmin = 0 rsw = 0 rswmin = 0
+ prwb = 0.1 prwg = 0.052 wr = 1
+ voff = -0.1819 voffl = 0 minv = 0
+ nfactor = 2.5373 eta0 = 0.2 etab = -2.5E-4
+ dsub = 1 cit = -6.393105E-11 cdsc = 2.8125E-7
+ cdscb = 1E-4 cdscd = 1E-10 pclm = 0.030097
+ pdiblc1 = 0 pdiblc2 = 2.76795476116616E-3 lpdiblc2 = -7.918431740325089E-10
+ wpdiblc2 = -4.490334098597363E-9 ppdiblc2 = 2.584364367796898E-14 pdiblcb = -0.025
+ drout = 0.43496 pscbe1 = 8E8 pscbe2 = 8.6797E-9
+ pvag = 0 delta = 0.019014310076038 ldelta = 4.376675112517461E-8
+ wdelta = -1.560184732591747E-8 pdelta = 3.352079855773622E-14 fprout = 0
+ pdits = 0 pditsl = 0 pditsd = 0
+ lambda = 0 vtl = 0 lc = 5E-9
+ xn = 3 alpha0 = 5.0449517E-13 alpha1 = -4.0583656E-18
+ beta0 = 6.2016506 aigbacc = 0.43 bigbacc = 0.054
+ cigbacc = 0.075 nigbacc = 1 aigbinv = 0.35
+ bigbinv = 0.03 cigbinv = 6E-3 eigbinv = 1.1
+ nigbinv = 3 aigc = 0.43 bigc = 0.054
+ cigc = 0.075 aigsd = 0.43 bigsd = 0.054
+ cigsd = 0.075 dlcig = 0 nigc = 1
+ poxedge = 1 pigcd = 1 ntox = 1
+ toxref = 4.23E-9 agidl = 0 bgidl = 2.3E9
+ cgidl = 0.5 egidl = 0.8 noia = 3E41
+ noib = 0 noic = 0 em = 4.1E7
+ af = 1 ef = 0.88 kf = 0
+ lintnoi = 0 tnoia = 2.5E7 tnoib = 0
+ ntnoi = 1 rnoia = 0.69 rnoib = 0.34
+ xpart = 0 cgso = {2E-11/sw_func_tox_lv_ratio} cgdo = {2E-11/sw_func_tox_lv_ratio}
+ cgbo = {1E-13/sw_func_tox_lv_ratio} ckappas = 0.6 cf = 0
+ clc = 7E-8 cle = 0.492 dlc = -1.2E-8
+ dwc = 0 vfbcv = -1 noff = 2.6123
+ voffcv = 0.112 acde = 0.44 moin = 8.7
+ cgsl = {0/sw_func_tox_lv_ratio} cgdl = {0/sw_func_tox_lv_ratio} ijthsrev = 0.1
+ ijthsfwd = 0.1 xjbvs = 1 bvs = 12.69
+ jss = 2.1483E-5 jsws = 1.4472E-10 cjs = {7.682E-04*sw_func_psd_nw_cj}
+ mjs = 0.3362 mjsws = 0.2659 cjsws = {9.160236799999998E-11*sw_func_psd_nw_cj}
+ cjswgs = {2.39155046E-10*sw_func_psd_nw_cj} mjswgs = 0.9274 pbs = 0.6587
+ pbsws = 0.7418 pbswgs = 1.4338 xrcrg1 = 12
+ xrcrg2 = 1 rbpb = 50 rbpd = 50
+ rbps = 50 rbdb = 50 rbsb = 50
+ gbmin = 1E-12 tnom = 30 ute = -0.450297722
+ lute = 1.2674939087568E-6 kt1 = -0.591648830672 lkt1 = 1.193649236237272E-9
+ wkt1 = -5.876714542820746E-8 pkt1 = 2.347394856984318E-13 kt1l = 0
+ kt2 = -0.055045 ua1 = 6.68269488E-10 lua1 = 1.111262531327999E-16
+ ub1 = -1.537629898795256E-19 lub1 = 2.904357429287962E-26 wub1 = -7.336489817770183E-26
+ pub1 = 5.865083419918195E-31 uc1 = -9.961E-12 at = 3.018023377950719E5
+ lat = -0.119002514088636 wat = -0.02491726966156 pat = 9.952954193613557E-8
+ prt = 0 njs = 1.3632 xtis = 5.2
+ tpb = 1.671E-3 tpbsw = 1.246E-3 tpbswg = 0
+ tcj = 1.2407E-3 tcjsw = 3.7357E-4 tcjswg = 2E-12
+ tvoff = 0 tvfbsdoff = 0 saref = 3E-6
+ sbref = 3E-6 wlod = 0 ku0 = 5.9E-8
+ kvsat = 0 kvth0 = 1.76E-8 tku0 = 0
+ llodku0 = 0 wlodku0 = 1 llodvth = 0
+ wlodvth = 1 lku0 = 0 wku0 = 0
+ pku0 = 0 lkvth0 = 0 wkvth0 = 7.3E-7
+ pkvth0 = 0 stk2 = 0 lodk2 = 1
+ steta0 = 0 lodeta0 = 1

.model plowvt_model.24 pmos
+ level = 54 lmin = 2E-6 lmax = 4E-6 wmin = 1E-6
+ wmax = 3E-6 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 4.23E-9
+ toxm = 4.23E-9 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 9.999999999999999E22 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {7.476E-9+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {2.8E-9-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = -7.916E-9 dwb = 0 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = -0.44077853074449 lvth0 = 4.524815608631753E-8
+ wvth0 = 5.395326185049154E-8 pvth0 = -5.874543012458974E-14 k1 = 0.64774
+ k2 = -0.042154641543781 lk2 = -1.418978714070311E-8 wk2 = 9.740546259168554E-9
+ pk2 = -4.903534003850292E-15 k3 = 3.39 k3b = 1
+ w0 = 1E-8 lpe0 = 0 lpeb = 0
+ vbm = -3 dvtp0 = 0 dvtp1 = 0
+ dvt0 = 2.4422 dvt1 = 0.16136 dvt2 = 0.026237
+ dvt0w = 0.5 dvt1w = 1.9281E6 dvt2w = -0.032
+ vfbsdoff = 0 u0 = 2.687485181380054E-3 lu0 = -2.379421229037608E-10
+ wu0 = -2.259049024626954E-10 pu0 = 6.523639197937554E-16 ua = -2.84069861096E-9
+ lua = -9.809146597881605E-17 wua = -1.432864503510736E-16 pua = 2.928077343371329E-22
+ ub = 2.8031381739656E-18 lub = 1.186906738343677E-25 wub = 2.760029888803342E-25
+ pub = -3.542973585479316E-31 uc = 7.363920700586722E-11 luc = -5.79582437008696E-17
+ wuc = -8.917843454715497E-18 puc = 5.709165204105419E-23 ud = 0
+ up = 0 lp = 1 eu = 1.67
+ vsat = 1.2376E5 a0 = 2.173045337634465 la0 = -1.08866813456044E-6
+ wa0 = -4.85276840350078E-7 pa0 = 6.302803604700511E-13 ags = 0.438644385795122
+ lags = -2.93628162139826E-8 wags = -1.732552957284442E-7 pags = 2.71708009000799E-13
+ b0 = 0 b1 = 2.1073E-24 keta = -0.01258
+ a1 = 0 a2 = 0.46703705 rdsw = 484.7
+ rdswmin = 0 rdw = 0 rdwmin = 0
+ rsw = 0 rswmin = 0 prwb = 0.1
+ prwg = 0.052 wr = 1 voff = -0.1819
+ voffl = 0 minv = 0 nfactor = 2.5373
+ eta0 = 0.2 etab = -2.5E-4 dsub = 1
+ cit = -6.393105E-11 cdsc = 2.8125E-7 cdscb = 1E-4
+ cdscd = 1E-10 pclm = 0.030097 pdiblc1 = 0
+ pdiblc2 = 7.195206015199029E-6 lpdiblc2 = 1.023573479306249E-8 wpdiblc2 = 5.542977376499927E-12
+ ppdiblc2 = 7.88531228569898E-15 pdiblcb = -0.025 drout = 0.43496
+ pscbe1 = 8E8 pscbe2 = 8.6797E-9 pvag = 0
+ delta = 0.012139940837888 ldelta = 7.122573161004257E-8 wdelta = 8.975747882217698E-9
+ pdelta = -6.465194774163889E-14 fprout = 0 pdits = 0
+ pditsl = 0 pditsd = 0 lambda = 0
+ vtl = 0 lc = 5E-9 xn = 3
+ alpha0 = 5.0449517E-13 alpha1 = -4.0583656E-18 beta0 = 6.2016506
+ aigbacc = 0.43 bigbacc = 0.054 cigbacc = 0.075
+ nigbacc = 1 aigbinv = 0.35 bigbinv = 0.03
+ cigbinv = 6E-3 eigbinv = 1.1 nigbinv = 3
+ aigc = 0.43 bigc = 0.054 cigc = 0.075
+ aigsd = 0.43 bigsd = 0.054 cigsd = 0.075
+ dlcig = 0 nigc = 1 poxedge = 1
+ pigcd = 1 ntox = 1 toxref = 4.23E-9
+ agidl = 0 bgidl = 2.3E9 cgidl = 0.5
+ egidl = 0.8 noia = 3E41 noib = 0
+ noic = 0 em = 4.1E7 af = 1
+ ef = 0.88 kf = 0 lintnoi = 0
+ tnoia = 2.5E7 tnoib = 0 ntnoi = 1
+ rnoia = 0.69 rnoib = 0.34 xpart = 0
+ cgso = {2E-11/sw_func_tox_lv_ratio} cgdo = {2E-11/sw_func_tox_lv_ratio} cgbo = {1E-13/sw_func_tox_lv_ratio}
+ ckappas = 0.6 cf = 0 clc = 7E-8
+ cle = 0.492 dlc = -1.2E-8 dwc = 0
+ vfbcv = -1 noff = 2.6123 voffcv = 0.112
+ acde = 0.44 moin = 8.7 cgsl = {0/sw_func_tox_lv_ratio}
+ cgdl = {0/sw_func_tox_lv_ratio} ijthsrev = 0.1 ijthsfwd = 0.1
+ xjbvs = 1 bvs = 12.69 jss = 2.1483E-5
+ jsws = 1.4472E-10 cjs = {7.682E-04*sw_func_psd_nw_cj} mjs = 0.3362
+ mjsws = 0.2659 cjsws = {9.160236799999998E-11*sw_func_psd_nw_cj} cjswgs = {2.39155046E-10*sw_func_psd_nw_cj}
+ mjswgs = 0.9274 pbs = 0.6587 pbsws = 0.7418
+ pbswgs = 1.4338 xrcrg1 = 12 xrcrg2 = 1
+ rbpb = 50 rbpd = 50 rbps = 50
+ rbdb = 50 rbsb = 50 gbmin = 1E-12
+ tnom = 30 ute = -0.143431564169984 lute = 4.174772792058415E-8
+ wute = 3.119842072248243E-8 pute = -1.246189717338838E-13 kt1 = -0.59135
+ kt1l = 0 kt2 = -0.055045 ua1 = 6.9609E-10
+ ub1 = -1.710349202409488E-19 lub1 = 9.803457292854824E-26 wub1 = 1.467297963554037E-25
+ pub1 = -2.926379058512171E-31 uc1 = -9.961E-12 at = 3.03830652E5
+ lat = -0.1271044123488 prt = 0 njs = 1.3632
+ xtis = 5.2 tpb = 1.671E-3 tpbsw = 1.246E-3
+ tpbswg = 0 tcj = 1.2407E-3 tcjsw = 3.7357E-4
+ tcjswg = 2E-12 tvoff = 0 tvfbsdoff = 0
+ saref = 3E-6 sbref = 3E-6 wlod = 0
+ ku0 = 5.9E-8 kvsat = 0 kvth0 = 1.76E-8
+ tku0 = 0 llodku0 = 0 wlodku0 = 1
+ llodvth = 0 wlodvth = 1 lku0 = 0
+ wku0 = 0 pku0 = 0 lkvth0 = 0
+ wkvth0 = 7.3E-7 pkvth0 = 0 stk2 = 0
+ lodk2 = 1 steta0 = 0 lodeta0 = 1

.model plowvt_model.25 pmos
+ level = 54 lmin = 1.5E-6 lmax = 2E-6 wmin = 1E-6
+ wmax = 3E-6 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 4.23E-9
+ toxm = 4.23E-9 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 9.999999999999999E22 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {7.476E-9+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {2.8E-9-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = -7.916E-9 dwb = 0 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = -0.340457164511725 lvth0 = -1.548327767283086E-7
+ wvth0 = -1.336740037016543E-7 pvth0 = 3.1545838829261E-13 k1 = 0.64774
+ k2 = -0.022732358293777 lk2 = -5.292558885451132E-8 wk2 = -4.066112633301831E-8
+ pk2 = 9.561756181400718E-14 k3 = 3.39 k3b = 1
+ w0 = 1E-8 lpe0 = 0 lpeb = 0
+ vbm = -3 dvtp0 = 0 dvtp1 = 0
+ dvt0 = 2.4422 dvt1 = 0.16136 dvt2 = 0.026237
+ dvt0w = 0.5 dvt1w = 1.9281E6 dvt2w = -0.032
+ vfbsdoff = 0 u0 = 2.442512659830791E-3 lu0 = 2.506310740740881E-10
+ wu0 = 2.233856496783778E-10 pu0 = -2.43701157396401E-16 ua = -2.8863E-9
+ ub = 2.8626501444E-18 wub = 9.835690055906879E-26 uc = 4.457871578E-11
+ wuc = 1.970813530634255E-17 ud = 0 up = 0
+ lp = 1 eu = 1.67 vsat = 1.2376E5
+ a0 = 1.96540299396057 la0 = -6.745462443372222E-7 wa0 = -2.982554516587431E-7
+ pa0 = 2.572849028640529E-13 ags = 0.219550011043712 lags = 4.075990047902291E-7
+ wags = 3.104566025318987E-8 pags = -1.357498176089718E-13 b0 = 0
+ b1 = 2.1073E-24 keta = -0.01258 a1 = 0
+ a2 = 0.46703705 rdsw = 484.7 rdswmin = 0
+ rdw = 0 rdwmin = 0 rsw = 0
+ rswmin = 0 prwb = 0.1 prwg = 0.052
+ wr = 1 voff = -0.1819 voffl = 0
+ minv = 0 nfactor = 2.5373 eta0 = 0.2
+ etab = -2.5E-4 dsub = 1 cit = -6.393105E-11
+ cdsc = 2.8125E-7 cdscb = 1E-4 cdscd = 1E-10
+ pclm = 0.030097 pdiblc1 = 0 pdiblc2 = 0.010890299145371
+ lpdiblc2 = -1.146952770358847E-8 wpdiblc2 = -2.705205417224337E-8 ppdiblc2 = 6.184898404090085E-14
+ pdiblcb = -0.025 drout = 0.43496 pscbe1 = 8E8
+ pscbe2 = 8.6797E-9 pvag = 0 delta = 0.101633746222899
+ ldelta = -1.072607138498237E-7 wdelta = -1.432520780693168E-7 pdelta = 2.389512283361015E-13
+ fprout = 0 pdits = 0 pditsl = 0
+ pditsd = 0 lambda = 0 vtl = 0
+ lc = 5E-9 xn = 3 alpha0 = 5.0449517E-13
+ alpha1 = -4.0583656E-18 beta0 = 6.2016506 aigbacc = 0.43
+ bigbacc = 0.054 cigbacc = 0.075 nigbacc = 1
+ aigbinv = 0.35 bigbinv = 0.03 cigbinv = 6E-3
+ eigbinv = 1.1 nigbinv = 3 aigc = 0.43
+ bigc = 0.054 cigc = 0.075 aigsd = 0.43
+ bigsd = 0.054 cigsd = 0.075 dlcig = 0
+ nigc = 1 poxedge = 1 pigcd = 1
+ ntox = 1 toxref = 4.23E-9 agidl = 0
+ bgidl = 2.3E9 cgidl = 0.5 egidl = 0.8
+ noia = 3E41 noib = 0 noic = 0
+ em = 4.1E7 af = 1 ef = 0.88
+ kf = 0 lintnoi = 0 tnoia = 2.5E7
+ tnoib = 0 ntnoi = 1 rnoia = 0.69
+ rnoib = 0.34 xpart = 0 cgso = {2E-11/sw_func_tox_lv_ratio}
+ cgdo = {2E-11/sw_func_tox_lv_ratio} cgbo = {1E-13/sw_func_tox_lv_ratio} ckappas = 0.6
+ cf = 0 clc = 7E-8 cle = 0.492
+ dlc = -1.2E-8 dwc = 0 vfbcv = -1
+ noff = 2.6123 voffcv = 0.112 acde = 0.44
+ moin = 8.7 cgsl = {0/sw_func_tox_lv_ratio} cgdl = {0/sw_func_tox_lv_ratio}
+ ijthsrev = 0.1 ijthsfwd = 0.1 xjbvs = 1
+ bvs = 12.69 jss = 2.1483E-5 jsws = 1.4472E-10
+ cjs = {7.682E-04*sw_func_psd_nw_cj} mjs = 0.3362 mjsws = 0.2659
+ cjsws = {9.160236799999998E-11*sw_func_psd_nw_cj} cjswgs = {2.39155046E-10*sw_func_psd_nw_cj} mjswgs = 0.9274
+ pbs = 0.6587 pbsws = 0.7418 pbswgs = 1.4338
+ xrcrg1 = 12 xrcrg2 = 1 rbpb = 50
+ rbpd = 50 rbps = 50 rbdb = 50
+ rbsb = 50 gbmin = 1E-12 tnom = 30
+ ute = -0.129255825086208 lute = 1.347563389190118E-8 wute = -1.111684087806509E-8
+ pute = -4.022541399775184E-14 kt1 = -0.629505684552704 lkt1 = 7.609769727191266E-8
+ wkt1 = 1.138965498626797E-7 pkt1 = -2.271552790461284E-13 kt1l = 0
+ kt2 = -0.026684374282701 lkt2 = -5.656243193058148E-8 wkt2 = -8.465782907617251E-8
+ pkt2 = 1.688415743095185E-13 ua1 = 6.15656874847232E-10 lua1 = 1.604158248046805E-16
+ wua1 = 2.400967393710199E-16 pua1 = -4.788489370015621E-22 ub1 = 4.142986281932788E-20
+ lub1 = -3.257051904068676E-25 wub1 = -4.874877793891093E-25 pub1 = 9.722456272136397E-31
+ uc1 = -9.961E-12 at = 2.250791940567041E5 lat = 0.029957495373309
+ wat = 0.237636011441888 pat = -4.73941261219701E-7 prt = 0
+ njs = 1.3632 xtis = 5.2 tpb = 1.671E-3
+ tpbsw = 1.246E-3 tpbswg = 0 tcj = 1.2407E-3
+ tcjsw = 3.7357E-4 tcjswg = 2E-12 tvoff = 0
+ tvfbsdoff = 0 saref = 3E-6 sbref = 3E-6
+ wlod = 0 ku0 = 5.9E-8 kvsat = 0
+ kvth0 = 1.76E-8 tku0 = 0 llodku0 = 0
+ wlodku0 = 1 llodvth = 0 wlodvth = 1
+ lku0 = 0 wku0 = 0 pku0 = 0
+ lkvth0 = 0 wkvth0 = 7.3E-7 pkvth0 = 0
+ stk2 = 0 lodk2 = 1 steta0 = 0
+ lodeta0 = 1

.model plowvt_model.26 pmos
+ level = 54 lmin = 1E-6 lmax = 1.5E-6 wmin = 1E-6
+ wmax = 3E-6 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 4.23E-9
+ toxm = 4.23E-9 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 9.999999999999999E22 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {7.476E-9+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {2.8E-9-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = -7.916E-9 dwb = 0 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = -0.405183643969011 lvth0 = -5.810552582733995E-8
+ wvth0 = 3.911886051638663E-8 pvth0 = 5.723673200516955E-14 k1 = 0.64774
+ k2 = -0.067353100424851 lk2 = 1.375564818616547E-8 wk2 = 3.238995473529882E-8
+ pk2 = -1.354997373448592E-14 k3 = 3.39 k3b = 1
+ w0 = 1E-8 lpe0 = 0 lpeb = 0
+ vbm = -3 dvtp0 = 0 dvtp1 = 0
+ dvt0 = 2.4422 dvt1 = 0.16136 dvt2 = 0.026237
+ dvt0w = 0.5 dvt1w = 1.9281E6 dvt2w = -0.032
+ vfbsdoff = 0 u0 = 4.492034960573883E-4 lu0 = 3.229432288417061E-9
+ wu0 = 2.189020459263662E-9 pu0 = -3.181145816840649E-15 ua = -3.20660305331904E-9
+ lua = 4.733078560025336E-16 wua = 3.155138820658143E-16 pua = -4.662309569395837E-22
+ ub = 2.75549336890368E-18 lub = 1.601350853017012E-25 wub = 2.039114679481682E-25
+ pub = -1.577407455062702E-31 uc = -5.239965021003523E-11 luc = 1.449244701355086E-16
+ wuc = 1.152364807680948E-16 puc = -1.427575594580425E-22 ud = 0
+ up = 0 lp = 1 eu = 1.67
+ vsat = 1.2376E5 a0 = 1.96466058591586 la0 = -6.73436789755208E-7
+ wa0 = -5.699917070192458E-7 pa0 = 6.633675628747881E-13 ags = 0.302208987013952
+ lags = 2.840734311003019E-7 wags = 1.274563585598804E-7 pags = -2.798259651584901E-13
+ b0 = 0 b1 = 2.1073E-24 keta = -0.01258
+ a1 = 0 a2 = 0.46703705 rdsw = 484.7
+ rdswmin = 0 rdw = 0 rdwmin = 0
+ rsw = 0 rswmin = 0 prwb = 0.1
+ prwg = 0.052 wr = 1 voff = -0.1819
+ voffl = 0 minv = 0 nfactor = -1.69910304676864
+ lnfactor = 6.330880713091056E-6 wnfactor = 4.173060348413355E-6 pnfactor = -6.236221384668918E-12
+ eta0 = 0.2 etab = -2.5E-4 dsub = 1
+ cit = -6.393105E-11 cdsc = 2.8125E-7 cdscb = 1E-4
+ cdscd = 1E-10 pclm = 0.030097 pdiblc1 = 0
+ pdiblc2 = -9.220234964289283E-3 lpdiblc2 = 1.858365446988767E-8 wpdiblc2 = 2.658470687510323E-8
+ ppdiblc2 = -1.83057916682539E-14 pdiblcb = -0.025 drout = 0.43496
+ pscbe1 = 8E8 pscbe2 = 8.6797E-9 pvag = 0
+ delta = -0.030526129135802 ldelta = 9.023900388621872E-8 wdelta = 7.612759178896309E-8
+ pdelta = -8.888975030011197E-14 fprout = 0 pdits = 0
+ pditsl = 0 pditsd = 0 lambda = 0
+ vtl = 0 lc = 5E-9 xn = 3
+ alpha0 = 5.0449517E-13 alpha1 = -4.0583656E-18 beta0 = 6.2016506
+ aigbacc = 0.43 bigbacc = 0.054 cigbacc = 0.075
+ nigbacc = 1 aigbinv = 0.35 bigbinv = 0.03
+ cigbinv = 6E-3 eigbinv = 1.1 nigbinv = 3
+ aigc = 0.43 bigc = 0.054 cigc = 0.075
+ aigsd = 0.43 bigsd = 0.054 cigsd = 0.075
+ dlcig = 0 nigc = 1 poxedge = 1
+ pigcd = 1 ntox = 1 toxref = 4.23E-9
+ agidl = 0 bgidl = 2.3E9 cgidl = 0.5
+ egidl = 0.8 noia = 3E41 noib = 0
+ noic = 0 em = 4.1E7 af = 1
+ ef = 0.88 kf = 0 lintnoi = 0
+ tnoia = 2.5E7 tnoib = 0 ntnoi = 1
+ rnoia = 0.69 rnoib = 0.34 xpart = 0
+ cgso = {2E-11/sw_func_tox_lv_ratio} cgdo = {2E-11/sw_func_tox_lv_ratio} cgbo = {1E-13/sw_func_tox_lv_ratio}
+ ckappas = 0.6 cf = 0 clc = 7E-8
+ cle = 0.492 dlc = -1.2E-8 dwc = 0
+ vfbcv = -1 noff = 2.6123 voffcv = 0.112
+ acde = 0.44 moin = 8.7 cgsl = {0/sw_func_tox_lv_ratio}
+ cgdl = {0/sw_func_tox_lv_ratio} ijthsrev = 0.1 ijthsfwd = 0.1
+ xjbvs = 1 bvs = 12.69 jss = 2.1483E-5
+ jsws = 1.4472E-10 cjs = {7.682E-04*sw_func_psd_nw_cj} mjs = 0.3362
+ mjsws = 0.2659 cjsws = {9.160236799999998E-11*sw_func_psd_nw_cj} cjswgs = {2.39155046E-10*sw_func_psd_nw_cj}
+ mjswgs = 0.9274 pbs = 0.6587 pbsws = 0.7418
+ pbswgs = 1.4338 xrcrg1 = 12 xrcrg2 = 1
+ rbpb = 50 rbpd = 50 rbps = 50
+ rbdb = 50 rbsb = 50 gbmin = 1E-12
+ tnom = 30 ute = 0.600531906849984 lute = -1.077119152713544E-6
+ wute = -7.480276285787632E-7 pute = 1.061014067142171E-12 kt1 = -0.489533825984
+ lkt1 = -1.33076248173158E-7 wkt1 = -1.258262627421124E-7 pkt1 = 1.31086492110473E-13
+ kt1l = 0 kt2 = -0.121721846517299 lkt2 = 8.546156657680233E-8
+ wkt2 = 8.465782907617253E-8 pkt2 = -8.418374523334597E-14 ua1 = 8.851911571527682E-10
+ lua1 = -2.423762066727126E-16 wua1 = -2.4009673937102E-16 pua1 = 2.387521976305422E-22
+ ub1 = -5.05827334819328E-19 lub1 = 4.921159657443398E-25 wub1 = 4.874877793891093E-25
+ pub1 = -4.847578478245304E-31 uc1 = -9.961E-12 at = 3.41329329328192E5
+ lat = -0.143766706776402 wat = -0.174274031516077 pat = 1.416171069766814E-7
+ prt = 0 njs = 1.3632 xtis = 5.2
+ tpb = 1.671E-3 tpbsw = 1.246E-3 tpbswg = 0
+ tcj = 1.2407E-3 tcjsw = 3.7357E-4 tcjswg = 2E-12
+ tvoff = 0 tvfbsdoff = 0 saref = 2.74E-6
+ sbref = 2.74E-6 wlod = 0 ku0 = 5.9E-8
+ kvsat = 0 kvth0 = 1.76E-8 tku0 = 0
+ llodku0 = 0 wlodku0 = 1 llodvth = 0
+ wlodvth = 1 lku0 = 0 wku0 = 0
+ pku0 = 0 lkvth0 = 0 wkvth0 = 7.3E-7
+ pkvth0 = 0 stk2 = 0 lodk2 = 1
+ steta0 = 0 lodeta0 = 1

.model plowvt_model.27 pmos
+ level = 54 lmin = 5E-7 lmax = 1E-6 wmin = 1E-6
+ wmax = 3E-6 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 4.23E-9
+ toxm = 4.23E-9 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 9.999999999999999E22 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {7.476E-9+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {2.8E-9-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = -7.916E-9 dwb = 0 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = -0.478072690733466 lvth0 = 1.437534227523333E-8
+ wvth0 = 1.051285223451131E-7 pvth0 = -8.40327571731607E-15 k1 = 0.64774
+ k2 = -0.052382114766565 lk2 = -1.131499952434073E-9 wk2 = 1.99975950364738E-8
+ pk2 = -1.22701124997433E-15 k3 = 3.39 k3b = 1
+ w0 = 1E-8 lpe0 = 0 lpeb = 0
+ vbm = -3 dvtp0 = 0 dvtp1 = 0
+ dvt0 = 2.4422 dvt1 = 0.16136 dvt2 = 0.026237
+ dvt0w = 0.5 dvt1w = 1.9281E6 dvt2w = -0.032
+ vfbsdoff = 0 u0 = 4.002733598245011E-3 lu0 = -3.041980451983112E-10
+ wu0 = -1.26629982523618E-9 pu0 = 2.548246740659932E-16 ua = -2.705835824112001E-9
+ lua = -2.465507672094661E-17 wua = -1.388052570341214E-16 pua = -1.445600501860765E-23
+ ub = 2.955490879296E-18 lub = -3.874243903242257E-26 wub = -7.101691666076689E-26
+ pub = 1.156480401488549E-31 uc = 1.177368754403456E-10 luc = -2.425929097123007E-17
+ wuc = -4.480754371716156E-17 puc = 1.63902184900964E-23 ud = 0
+ up = 0 lp = 1 eu = 1.67
+ vsat = 1.238143166168397E5 lvsat = -5.40124437853698E-5 wvsat = 0.018634930202284
+ pvsat = -1.853057459315132E-8 a0 = 0.807693038289209 la0 = 4.770517396047334E-7
+ wa0 = 7.871910728520717E-7 pa0 = -6.862149934292501E-13 ags = 0.842872017209024
+ lags = -2.535618861256774E-7 wags = -2.350206176541785E-7 pags = 8.06211399887701E-14
+ b0 = 1.56750654074496E-6 lb0 = -1.558728504116788E-12 wb0 = -1.436732678991261E-12
+ pb0 = 1.42868697598891E-18 b1 = 5.445233442547199E-8 lb1 = -5.414740135268936E-14
+ wb1 = -1.625428319720863E-13 pb1 = 1.616325921130426E-19 keta = -0.01258
+ a1 = 0 a2 = 0.46703705 rdsw = 484.7
+ rdswmin = 0 rdw = 0 rdwmin = 0
+ rsw = 0 rswmin = 0 prwb = 0.1
+ prwg = 0.052 wr = 1 voff = -0.1819
+ voffl = 0 minv = 0 nfactor = 4.667430252799999
+ wnfactor = -2.098280545260134E-6 eta0 = 0.2 etab = -2.5E-4
+ dsub = 1 cit = -6.393105E-11 cdsc = 2.8125E-7
+ cdscb = 1E-4 cdscd = 1E-10 pclm = 0.030097
+ pdiblc1 = 0 pdiblc2 = -0.021380410164294 lpdiblc2 = 3.067573268877275E-8
+ wpdiblc2 = 7.611773786833068E-9 ppdiblc2 = 5.608929947219431E-16 pdiblcb = -0.025
+ drout = 0.43496 pscbe1 = 8E8 pscbe2 = 8.6797E-9
+ pvag = 0 delta = 0.051883719215571 ldelta = 8.290650685613601E-9
+ wdelta = -1.973334760553997E-8 pdelta = 6.434367833781882E-15 fprout = 0
+ pdits = 0 pditsl = 0 pditsd = 0
+ lambda = 0 vtl = 0 lc = 5E-9
+ xn = 3 alpha0 = 5.0449517E-13 alpha1 = -4.0583656E-18
+ beta0 = 6.2016506 aigbacc = 0.43 bigbacc = 0.054
+ cigbacc = 0.075 nigbacc = 1 aigbinv = 0.35
+ bigbinv = 0.03 cigbinv = 6E-3 eigbinv = 1.1
+ nigbinv = 3 aigc = 0.43 bigc = 0.054
+ cigc = 0.075 aigsd = 0.43 bigsd = 0.054
+ cigsd = 0.075 dlcig = 0 nigc = 1
+ poxedge = 1 pigcd = 1 ntox = 1
+ toxref = 4.23E-9 agidl = 0 bgidl = 2.3E9
+ cgidl = 0.5 egidl = 0.8 noia = 3E41
+ noib = 0 noic = 0 em = 4.1E7
+ af = 1 ef = 0.88 kf = 0
+ lintnoi = 0 tnoia = 2.5E7 tnoib = 0
+ ntnoi = 1 rnoia = 0.69 rnoib = 0.34
+ xpart = 0 cgso = {2E-11/sw_func_tox_lv_ratio} cgdo = {2E-11/sw_func_tox_lv_ratio}
+ cgbo = {1E-13/sw_func_tox_lv_ratio} ckappas = 0.6 cf = 0
+ clc = 7E-8 cle = 0.492 dlc = -1.2E-8
+ dwc = 0 vfbcv = -1 noff = 2.6123
+ voffcv = 0.112 acde = 0.44 moin = 8.7
+ cgsl = {0/sw_func_tox_lv_ratio} cgdl = {0/sw_func_tox_lv_ratio} ijthsrev = 0.1
+ ijthsfwd = 0.1 xjbvs = 1 bvs = 12.69
+ jss = 2.1483E-5 jsws = 1.4472E-10 cjs = {7.682E-04*sw_func_psd_nw_cj}
+ mjs = 0.3362 mjsws = 0.2659 cjsws = {9.160236799999998E-11*sw_func_psd_nw_cj}
+ cjswgs = {2.39155046E-10*sw_func_psd_nw_cj} mjswgs = 0.9274 pbs = 0.6587
+ pbsws = 0.7418 pbswgs = 1.4338 xrcrg1 = 12
+ xrcrg2 = 1 rbpb = 50 rbpd = 50
+ rbps = 50 rbdb = 50 rbsb = 50
+ gbmin = 1E-12 tnom = 30 ute = -0.43312091239008
+ lute = -4.925478926122441E-8 wute = 3.438932440570795E-7 pute = -2.47920486069107E-14
+ kt1 = -0.579089950839296 lkt1 = -4.402163761705209E-8 wkt1 = -1.714511620062926E-8
+ pkt1 = 2.301395998962209E-14 kt1l = 0 kt2 = -0.020754184
+ lkt2 = -1.49406770304E-8 ua1 = 3.8940488E-10 lua1 = 2.50633667328E-16
+ ub1 = 6.06298624E-19 lub1 = -6.137820877055999E-25 uc1 = -2.284941472E-11
+ luc1 = 1.2816239597568E-17 at = 3.280447318915072E5 lat = -0.130556503085363
+ wat = -0.060179739882998 pat = 2.816174337674791E-8 prt = 0
+ njs = 1.3632 xtis = 5.2 tpb = 1.671E-3
+ tpbsw = 1.246E-3 tpbswg = 0 tcj = 1.2407E-3
+ tcjsw = 3.7357E-4 tcjswg = 2E-12 tvoff = 0
+ tvfbsdoff = 0 saref = 2.74E-6 sbref = 2.74E-6
+ wlod = 0 ku0 = 5.9E-8 kvsat = 0
+ kvth0 = 1.76E-8 tku0 = 0 llodku0 = 0
+ wlodku0 = 1 llodvth = 0 wlodvth = 1
+ lku0 = 0 wku0 = 0 pku0 = 0
+ lkvth0 = 0 wkvth0 = 7.3E-7 pkvth0 = 0
+ stk2 = 0 lodk2 = 1 steta0 = 0
+ lodeta0 = 1

.model plowvt_model.28 pmos
+ level = 54 lmin = 3.5E-7 lmax = 5E-7 wmin = 1E-6
+ wmax = 3E-6 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 4.23E-9
+ toxm = 4.23E-9 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 9.999999999999999E22 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {7.476E-9+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {2.8E-9-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = -7.916E-9 dwb = 0 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = -0.545833552299904 lvth0 = 4.787631223368058E-8
+ wvth0 = 2.27209580137852E-7 pvth0 = -6.876015069004617E-14 k1 = 0.64774
+ k2 = -0.092880852834961 lk2 = 1.88910761485806E-8 wk2 = 3.475633437359948E-8
+ pk2 = -8.523731978249262E-15 k3 = 3.39 k3b = 1
+ w0 = 1E-8 lpe0 = 0 lpeb = 0
+ vbm = -3 dvtp0 = 0 dvtp1 = 0
+ dvt0 = 2.4422 dvt1 = 0.16136 dvt2 = 0.026237
+ dvt0w = 0.5 dvt1w = 1.9281E6 dvt2w = -0.032
+ vfbsdoff = 0 u0 = 3.487838784315712E-3 lu0 = -4.963404919166562E-11
+ wu0 = -1.345330519890127E-9 pu0 = 2.938974495029049E-16 ua = -2.321180996399998E-9
+ lua = -2.148284235417607E-16 wua = -5.056044559381749E-16 pua = 1.668895189195564E-22
+ ub = 2.016844243702399E-18 lub = 4.253244576050536E-25 wub = 5.068723631286392E-25
+ pub = -1.700604197790275E-31 uc = 1.17494276833792E-10 luc = -2.413935022014996E-17
+ wuc = -5.975131427857313E-17 puc = 2.377841865565828E-23 ud = 0
+ up = 0 lp = 1 eu = 1.67
+ vsat = 1.027510386533824E5 lvsat = 0.010359672181348 wvsat = 6.114509477842946E-3
+ pvsat = -1.234047858698761E-8 a0 = 2.037631514944256 la0 = -1.310298432535218E-7
+ wa0 = -8.618495389328095E-7 pa0 = 1.290706850371952E-13 ags = 0.33000412456
+ wags = -7.195196880957884E-8 b0 = -5.423438129831039E-6 lb0 = 1.897594541015986E-12
+ wb0 = 5.381391191087885E-12 pb0 = -1.94219346537822E-18 b1 = 5.127462474016005E-8
+ lb1 = -5.25763416842711E-14 wb1 = -1.530572160313651E-13 pb1 = 1.569429035919501E-19
+ keta = -0.01172621949648 lketa = -4.221090809402873E-10 wketa = -2.548575784471364E-9
+ pketa = 1.260015867842643E-15 a1 = 0 a2 = 0.46703705
+ rdsw = 484.7 rdswmin = 0 rdw = 0
+ rdwmin = 0 rsw = 0 rswmin = 0
+ prwb = 0.1 prwg = 0.052 wr = 1
+ voff = -0.1819 voffl = 0 minv = 0
+ nfactor = 4.667430252799999 wnfactor = -2.098280545260134E-6 eta0 = 0.2
+ etab = -2.5E-4 dsub = 1 cit = -6.393105E-11
+ cdsc = 2.8125E-7 cdscb = 1E-4 cdscd = 1E-10
+ pclm = 0.030097 pdiblc1 = 0 pdiblc2 = -0.096665417519808
+ lpdiblc2 = 6.789664032533866E-8 wpdiblc2 = 4.765677346437981E-8 ppdiblc2 = -1.923735484585716E-14
+ pdiblcb = -0.025 drout = 0.43496 pscbe1 = 8E8
+ pscbe2 = 8.6797E-9 pvag = 0 delta = -0.015351336128768
+ ldelta = 4.15316620478549E-8 wdelta = 9.840399425471464E-8 pdelta = -5.1972733981928E-14
+ fprout = 0 pdits = 0 pditsl = 0
+ pditsd = 0 lambda = 0 vtl = 0
+ lc = 5E-9 xn = 3 alpha0 = 5.0449517E-13
+ alpha1 = -4.0583656E-18 beta0 = 6.2016506 aigbacc = 0.43
+ bigbacc = 0.054 cigbacc = 0.075 nigbacc = 1
+ aigbinv = 0.35 bigbinv = 0.03 cigbinv = 6E-3
+ eigbinv = 1.1 nigbinv = 3 aigc = 0.43
+ bigc = 0.054 cigc = 0.075 aigsd = 0.43
+ bigsd = 0.054 cigsd = 0.075 dlcig = 0
+ nigc = 1 poxedge = 1 pigcd = 1
+ ntox = 1 toxref = 4.23E-9 agidl = 0
+ bgidl = 2.3E9 cgidl = 0.5 egidl = 0.8
+ noia = 3E41 noib = 0 noic = 0
+ em = 4.1E7 af = 1 ef = 0.88
+ kf = 0 lintnoi = 0 tnoia = 2.5E7
+ tnoib = 0 ntnoi = 1 rnoia = 0.69
+ rnoib = 0.34 xpart = 0 cgso = {2E-11/sw_func_tox_lv_ratio}
+ cgdo = {2E-11/sw_func_tox_lv_ratio} cgbo = {1E-13/sw_func_tox_lv_ratio} ckappas = 0.6
+ cf = 0 clc = 7E-8 cle = 0.492
+ dlc = -1.2E-8 dwc = 0 vfbcv = -1
+ noff = 2.6123 voffcv = 0.112 acde = 0.44
+ moin = 8.7 cgsl = {0/sw_func_tox_lv_ratio} cgdl = {0/sw_func_tox_lv_ratio}
+ ijthsrev = 0.1 ijthsfwd = 0.1 xjbvs = 1
+ bvs = 12.69 jss = 2.1483E-5 jsws = 1.4472E-10
+ cjs = {7.682E-04*sw_func_psd_nw_cj} mjs = 0.3362 mjsws = 0.2659
+ cjsws = {9.160236799999998E-11*sw_func_psd_nw_cj} cjswgs = {2.39155046E-10*sw_func_psd_nw_cj} mjswgs = 0.9274
+ pbs = 0.6587 pbsws = 0.7418 pbswgs = 1.4338
+ xrcrg1 = 12 xrcrg2 = 1 rbpb = 50
+ rbpd = 50 rbps = 50 rbdb = 50
+ rbsb = 50 gbmin = 1E-12 tnom = 30
+ ute = -0.63053937107168 lute = 4.83488967109586E-8 wute = 3.398919265598962E-7
+ pute = -2.281379723630328E-14 kt1 = -0.6776655255424 lkt1 = 4.714126516162574E-9
+ wkt1 = 1.45515285347302E-8 pkt1 = 7.343138832460378E-15 kt1l = 0
+ kt2 = -0.072560472589696 lkt2 = 1.06723520483457E-8 wkt2 = 9.898600834945484E-8
+ pkt2 = -4.893868252797048E-14 ua1 = 7.0051197668928E-10 lua1 = 9.682231872481998E-17
+ wua1 = 5.845858998076181E-16 pua1 = -2.890192688648864E-22 ub1 = -3.029774256080002E-19
+ lub1 = -1.642360087794048E-25 wub1 = -1.238000223781291E-24 pub1 = 6.120673106374701E-31
+ uc1 = 3.35229445113664E-11 luc1 = -1.505425480641955E-17 wuc1 = -9.089335194456524E-17
+ puc1 = 4.493767320139305E-23 at = 1.5108905364112E5 lat = -0.043069615758371
+ wat = -5.007351277669973E-3 pat = 8.845144502736446E-10 prt = 0
+ njs = 1.3632 xtis = 5.2 tpb = 1.671E-3
+ tpbsw = 1.246E-3 tpbswg = 0 tcj = 1.2407E-3
+ tcjsw = 3.7357E-4 tcjswg = 2E-12 tvoff = 0
+ tvfbsdoff = 0 saref = 1.74E-6 sbref = 1.74E-6
+ wlod = 0 ku0 = 5.9E-8 kvsat = 0
+ kvth0 = 1.76E-8 tku0 = 0 llodku0 = 0
+ wlodku0 = 1 llodvth = 0 wlodvth = 1
+ lku0 = 0 wku0 = 0 pku0 = 0
+ lkvth0 = 0 wkvth0 = 7.3E-7 pkvth0 = 0
+ stk2 = 0 lodk2 = 1 steta0 = 0
+ lodeta0 = 1

.model plowvt_model.29 pmos
+ level = 54 lmin = 8E-6 lmax = 2.02E-5 wmin = 5.5E-7
+ wmax = 1E-6 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 4.23E-9
+ toxm = 4.23E-9 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 9.999999999999999E22 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {7.476E-9+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {2.8E-9-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = -7.916E-9 dwb = 0 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = -0.434780795893333 wvth0 = 3.033336705713622E-8
+ k1 = 0.64774 k2 = -0.050907829104 wk2 = 1.206834424083699E-8
+ k3 = 3.39 k3b = 1 w0 = 1E-8
+ lpe0 = 0 lpeb = 0 vbm = -3
+ dvtp0 = 0 dvtp1 = 0 dvt0 = 2.4422
+ dvt1 = 0.16136 dvt2 = 0.026237 dvt0w = 0.5
+ dvt1w = 1.9281E6 dvt2w = -0.032 vfbsdoff = 0
+ u0 = 2.894566622862222E-3 wu0 = -3.323400479811863E-10 ua = -2.714727941333333E-9
+ wua = -1.690067132454827E-16 ub = 2.777107608888889E-18 wub = 1.604568240792175E-25
+ uc = 6.996144890666666E-11 wuc = -5.295075194614183E-18 ud = 0
+ up = 0 lp = 1 eu = 1.67
+ vsat = 1.2376E5 a0 = 1.177846302684444 wa0 = 2.921649386412935E-7
+ ags = 0.2878571328 wags = -1.243833191037436E-8 b0 = 9.975197112888891E-8
+ wb0 = -9.826047965656975E-14 b1 = -2.427691125333334E-7 wb1 = 2.391392287627349E-13
+ keta = -0.01258 a1 = 0 a2 = 0.46703705
+ rdsw = 484.7 rdswmin = 0 rdw = 0
+ rdwmin = 0 rsw = 0 rswmin = 0
+ prwb = 0.1 prwg = 0.052 wr = 1
+ voff = -0.1819 voffl = 0 minv = 0
+ nfactor = 2.5373 eta0 = 0.2 etab = -2.5E-4
+ dsub = 1 cit = -6.393105E-11 cdsc = 2.8125E-7
+ cdscb = 1E-4 cdscd = 1E-10 pclm = 0.030097
+ pdiblc1 = 0 pdiblc2 = 2.532779656533334E-3 wpdiblc2 = -1.123525709508847E-9
+ pdiblcb = -0.025 drout = 0.43496 pscbe1 = 8E8
+ pscbe2 = 8.6797E-9 pvag = 0 delta = 0.012113939964444
+ wdelta = 7.81202201903928E-10 fprout = 0 pdits = 0
+ pditsl = 0 pditsd = 0 lambda = 0
+ vtl = 0 lc = 5E-9 xn = 3
+ alpha0 = 5.0449517E-13 alpha1 = -4.0583656E-18 beta0 = 6.2016506
+ aigbacc = 0.43 bigbacc = 0.054 cigbacc = 0.075
+ nigbacc = 1 aigbinv = 0.35 bigbinv = 0.03
+ cigbinv = 6E-3 eigbinv = 1.1 nigbinv = 3
+ aigc = 0.43 bigc = 0.054 cigc = 0.075
+ aigsd = 0.43 bigsd = 0.054 cigsd = 0.075
+ dlcig = 0 nigc = 1 poxedge = 1
+ pigcd = 1 ntox = 1 toxref = 4.23E-9
+ agidl = 0 bgidl = 2.3E9 cgidl = 0.5
+ egidl = 0.8 noia = 3E41 noib = 0
+ noic = 0 em = 4.1E7 af = 1
+ ef = 0.88 kf = 0 lintnoi = 0
+ tnoia = 2.5E7 tnoib = 0 ntnoi = 1
+ rnoia = 0.69 rnoib = 0.34 xpart = 0
+ cgso = {2E-11/sw_func_tox_lv_ratio} cgdo = {2E-11/sw_func_tox_lv_ratio} cgbo = {1E-13/sw_func_tox_lv_ratio}
+ ckappas = 0.6 cf = 0 clc = 7E-8
+ cle = 0.492 dlc = -1.2E-8 dwc = 0
+ vfbcv = -1 noff = 2.6123 voffcv = 0.112
+ acde = 0.44 moin = 8.7 cgsl = {0/sw_func_tox_lv_ratio}
+ cgdl = {0/sw_func_tox_lv_ratio} ijthsrev = 0.1 ijthsfwd = 0.1
+ xjbvs = 1 bvs = 12.69 jss = 2.1483E-5
+ jsws = 1.4472E-10 cjs = {7.682E-04*sw_func_psd_nw_cj} mjs = 0.3362
+ mjsws = 0.2659 cjsws = {9.160236799999998E-11*sw_func_psd_nw_cj} cjswgs = {2.39155046E-10*sw_func_psd_nw_cj}
+ mjswgs = 0.9274 pbs = 0.6587 pbsws = 0.7418
+ pbswgs = 1.4338 xrcrg1 = 12 xrcrg2 = 1
+ rbpb = 50 rbpd = 50 rbps = 50
+ rbdb = 50 rbsb = 50 gbmin = 1E-12
+ tnom = 30 ute = -0.298681844088889 wute = 6.828199156071825E-9
+ kt1 = -0.558095436444444 wkt1 = -6.230878132127292E-8 kt1l = 0
+ kt2 = -0.055045 ua1 = 6.8217E-10 ub1 = -1.5013E-19
+ uc1 = -9.961E-12 at = 2.648074853333333E5 wat = 9.311180667370668E-3
+ prt = 0 njs = 1.3632 xtis = 5.2
+ tpb = 1.671E-3 tpbsw = 1.246E-3 tpbswg = 0
+ tcj = 1.2407E-3 tcjsw = 3.7357E-4 tcjswg = 2E-12
+ tvoff = 0 tvfbsdoff = 0 saref = 3E-6
+ sbref = 3E-6 wlod = 0 ku0 = 5.9E-8
+ kvsat = 0 kvth0 = 1.76E-8 tku0 = 0
+ llodku0 = 0 wlodku0 = 1 llodvth = 0
+ wlodvth = 1 lku0 = 0 wku0 = 0
+ pku0 = 0 lkvth0 = 0 wkvth0 = 7.3E-7
+ pkvth0 = 0 stk2 = 0 lodk2 = 1
+ steta0 = 0 lodeta0 = 1

.model plowvt_model.30 pmos
+ level = 54 lmin = 4E-6 lmax = 8E-6 wmin = 5.5E-7
+ wmax = 1E-6 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 4.23E-9
+ toxm = 4.23E-9 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 9.999999999999999E22 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {7.476E-9+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {2.8E-9-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = -7.916E-9 dwb = 0 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = -0.452351271317327 lvth0 = 1.404654087295738E-7
+ wvth0 = 3.349754334921872E-8 pvth0 = -2.529569094942426E-14 k1 = 0.64774
+ k2 = -0.051058193484518 lk2 = 1.202073003610587E-9 wk2 = 1.065104963347926E-8
+ pk2 = 1.133042000906067E-14 k3 = 3.39 k3b = 1
+ w0 = 1E-8 lpe0 = 0 lpeb = 0
+ vbm = -3 dvtp0 = 0 dvtp1 = 0
+ dvt0 = 2.4422 dvt1 = 0.16136 dvt2 = 0.026237
+ dvt0w = 0.5 dvt1w = 1.9281E6 dvt2w = -0.032
+ vfbsdoff = 0 u0 = 2.75321155871016E-3 lu0 = 1.130048924857243E-9
+ wu0 = -2.001799573955536E-10 pu0 = -1.056540628177782E-15 ua = -2.653280831004088E-9
+ lua = -4.912327788161127E-16 wua = -1.803516197410844E-16 pua = 9.069572048843802E-23
+ ub = 2.63224513268409E-18 lub = 1.158088579771648E-24 wub = 2.215087951174029E-25
+ pub = -4.880738772676691E-31 uc = 6.3542737727296E-11 luc = 5.131374465236087E-17
+ wuc = 1.027663415202534E-18 puc = -5.054650154231876E-23 ud = 0
+ up = 0 lp = 1 eu = 1.67
+ vsat = 1.2376E5 a0 = 0.932293362066481 la0 = 1.963048428476243E-6
+ wa0 = 4.419808615946533E-7 pa0 = -1.19768841445834E-12 ags = 0.148820416510155
+ lags = 1.11151512470754E-6 wags = 7.609053482896284E-8 pags = -7.077351722609573E-13
+ b0 = 2.33780943434951E-8 lb0 = 6.105633205731522E-13 wb0 = -2.302854507687117E-14
+ pb0 = -6.014341778039423E-19 b1 = -2.450250413607111E-7 lb1 = 1.803479741758876E-14
+ wb1 = 2.413614269422858E-13 pb1 = -1.776514112660097E-20 keta = -0.01258
+ a1 = 0 a2 = 0.46703705 rdsw = 484.7
+ rdswmin = 0 rdw = 0 rdwmin = 0
+ rsw = 0 rswmin = 0 prwb = 0.1
+ prwg = 0.052 wr = 1 voff = -0.1819
+ voffl = 0 minv = 0 nfactor = 2.5373
+ eta0 = 0.2 etab = -2.5E-4 dsub = 1
+ cit = -6.393105E-11 cdsc = 2.8125E-7 cdscb = 1E-4
+ cdscd = 1E-10 pclm = 0.030097 pdiblc1 = 0
+ pdiblc2 = -1.294702722331236E-3 lpdiblc2 = 3.059842512959491E-8 wpdiblc2 = -4.884214697932211E-10
+ ppdiblc2 = -5.077277333982598E-15 pdiblcb = -0.025 drout = 0.43496
+ pscbe1 = 8E8 pscbe2 = 8.6797E-9 pvag = 0
+ delta = -3.86990188027733E-3 ldelta = 1.277812252434438E-7 wdelta = 6.940199893227424E-9
+ pdelta = -4.923749114351655E-14 fprout = 0 pdits = 0
+ pditsl = 0 pditsd = 0 lambda = 0
+ vtl = 0 lc = 5E-9 xn = 3
+ alpha0 = 5.0449517E-13 alpha1 = -4.0583656E-18 beta0 = 6.2016506
+ aigbacc = 0.43 bigbacc = 0.054 cigbacc = 0.075
+ nigbacc = 1 aigbinv = 0.35 bigbinv = 0.03
+ cigbinv = 6E-3 eigbinv = 1.1 nigbinv = 3
+ aigc = 0.43 bigc = 0.054 cigc = 0.075
+ aigsd = 0.43 bigsd = 0.054 cigsd = 0.075
+ dlcig = 0 nigc = 1 poxedge = 1
+ pigcd = 1 ntox = 1 toxref = 4.23E-9
+ agidl = 0 bgidl = 2.3E9 cgidl = 0.5
+ egidl = 0.8 noia = 3E41 noib = 0
+ noic = 0 em = 4.1E7 af = 1
+ ef = 0.88 kf = 0 lintnoi = 0
+ tnoia = 2.5E7 tnoib = 0 ntnoi = 1
+ rnoia = 0.69 rnoib = 0.34 xpart = 0
+ cgso = {2E-11/sw_func_tox_lv_ratio} cgdo = {2E-11/sw_func_tox_lv_ratio} cgbo = {1E-13/sw_func_tox_lv_ratio}
+ ckappas = 0.6 cf = 0 clc = 7E-8
+ cle = 0.492 dlc = -1.2E-8 dwc = 0
+ vfbcv = -1 noff = 2.6123 voffcv = 0.112
+ acde = 0.44 moin = 8.7 cgsl = {0/sw_func_tox_lv_ratio}
+ cgdl = {0/sw_func_tox_lv_ratio} ijthsrev = 0.1 ijthsfwd = 0.1
+ xjbvs = 1 bvs = 12.69 jss = 2.1483E-5
+ jsws = 1.4472E-10 cjs = {7.682E-04*sw_func_psd_nw_cj} mjs = 0.3362
+ mjsws = 0.2659 cjsws = {9.160236799999998E-11*sw_func_psd_nw_cj} cjswgs = {2.39155046E-10*sw_func_psd_nw_cj}
+ mjswgs = 0.9274 pbs = 0.6587 pbsws = 0.7418
+ pbswgs = 1.4338 xrcrg1 = 12 xrcrg2 = 1
+ rbpb = 50 rbpd = 50 rbps = 50
+ rbdb = 50 rbsb = 50 gbmin = 1E-12
+ tnom = 30 ute = -0.41994262456522 lute = 9.69407183439978E-7
+ wute = -2.990122801793558E-8 pute = 2.936297325998848E-13 kt1 = -0.58807718306368
+ lkt1 = 2.396860751728152E-7 wkt1 = -6.228538976148828E-8 pkt1 = -1.870014855423186E-16
+ kt1l = 0 kt2 = -0.055045 ua1 = 6.68269488E-10
+ lua1 = 1.111262531327999E-16 ub1 = -2.875736060909972E-19 lub1 = 1.098779164533869E-24
+ wub1 = 5.844498170017593E-26 pub1 = -4.672325617038865E-31 uc1 = -9.961E-12
+ at = 2.543498940423112E5 lat = 0.083602167816948 wat = 0.02182566515221
+ pat = -1.000457947655958E-7 prt = 0 njs = 1.3632
+ xtis = 5.2 tpb = 1.671E-3 tpbsw = 1.246E-3
+ tpbswg = 0 tcj = 1.2407E-3 tcjsw = 3.7357E-4
+ tcjswg = 2E-12 tvoff = 0 tvfbsdoff = 0
+ saref = 3E-6 sbref = 3E-6 wlod = 0
+ ku0 = 5.9E-8 kvsat = 0 kvth0 = 1.76E-8
+ tku0 = 0 llodku0 = 0 wlodku0 = 1
+ llodvth = 0 wlodvth = 1 lku0 = 0
+ wku0 = 0 pku0 = 0 lkvth0 = 0
+ wkvth0 = 7.3E-7 pkvth0 = 0 stk2 = 0
+ lodk2 = 1 steta0 = 0 lodeta0 = 1

.model plowvt_model.31 pmos
+ level = 54 lmin = 2E-6 lmax = 4E-6 wmin = 5.5E-7
+ wmax = 1E-6 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 4.23E-9
+ toxm = 4.23E-9 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 9.999999999999999E22 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {7.476E-9+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {2.8E-9-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = -7.916E-9 dwb = 0 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = -0.39416526966205 lvth0 = -9.195275628226272E-8
+ wvth0 = 8.036962247756726E-9 pvth0 = 7.640405420225549E-14 k1 = 0.64774
+ k2 = -0.040365655487738 lk2 = -4.150820077072468E-8 wk2 = 7.978309122635443E-9
+ pk2 = 2.20064147055752E-14 k3 = 3.39 k3b = 1
+ w0 = 1E-8 lpe0 = 0 lpeb = 0
+ vbm = -3 dvtp0 = 0 dvtp1 = 0
+ dvt0 = 2.4422 dvt1 = 0.16136 dvt2 = 0.026237
+ dvt0w = 0.5 dvt1w = 1.9281E6 dvt2w = -0.032
+ vfbsdoff = 0 u0 = 2.84889857458337E-3 lu0 = 7.478367086532951E-10
+ wu0 = -3.849048426108357E-10 pu0 = -3.186755466738592E-16 ua = -2.897261180302223E-9
+ lua = 4.833223284203531E-16 wua = -8.75696045456563E-17 pua = -2.799127610081799E-22
+ ub = 3.077949919512889E-18 lub = -6.222346207373066E-25 wub = 5.300228552467881E-27
+ pub = 3.75549621019307E-31 uc = 7.638915888E-11 wuc = -1.162667804842624E-17
+ ud = 0 up = 0 lp = 1
+ eu = 1.67 vsat = 1.2376E5 a0 = 1.669704515991282
+ la0 = -9.824666847609807E-7 wa0 = 1.053802932789652E-8 pa0 = 5.256668347479932E-13
+ ags = 0.388022956950891 lags = 1.560444971710637E-7 wags = -1.233907584882922E-7
+ pags = 8.907290576548599E-14 b0 = 2.274418516783645E-7 lb0 = -2.045489517252501E-13
+ wb0 = -2.240411411120696E-13 pb0 = 2.014905357990542E-19 b1 = -2.396919111838579E-7
+ lb1 = -3.267857760833993E-15 wb1 = 2.361080377278368E-13 pb1 = 3.218996751594003E-21
+ keta = -0.01258 a1 = 0 a2 = 0.46703705
+ rdsw = 484.7 rdswmin = 0 rdw = 0
+ rdwmin = 0 rsw = 0 rswmin = 0
+ prwb = 0.1 prwg = 0.052 wr = 1
+ voff = -0.1819 voffl = 0 minv = 0
+ nfactor = 2.5373 eta0 = 0.2 etab = -2.5E-4
+ dsub = 1 cit = -6.393105E-11 cdsc = 2.8125E-7
+ cdscb = 1E-4 cdscd = 1E-10 pclm = 0.030097
+ pdiblc1 = 0 pdiblc2 = 1.212501190861511E-3 lpdiblc2 = 2.05836498187378E-8
+ wpdiblc2 = -1.18174127238439E-9 ppdiblc2 = -2.307880714512434E-15 pdiblcb = -0.025
+ drout = 0.43496 pscbe1 = 8E8 pscbe2 = 8.6797E-9
+ pvag = 0 delta = 0.03276109190496 ldelta = -1.853761633230821E-8
+ wdelta = -1.133707573409944E-8 pdelta = 2.376925862227785E-14 fprout = 0
+ pdits = 0 pditsl = 0 pditsd = 0
+ lambda = 0 vtl = 0 lc = 5E-9
+ xn = 3 alpha0 = 5.0449517E-13 alpha1 = -4.0583656E-18
+ beta0 = 6.2016506 aigbacc = 0.43 bigbacc = 0.054
+ cigbacc = 0.075 nigbacc = 1 aigbinv = 0.35
+ bigbinv = 0.03 cigbinv = 6E-3 eigbinv = 1.1
+ nigbinv = 3 aigc = 0.43 bigc = 0.054
+ cigc = 0.075 aigsd = 0.43 bigsd = 0.054
+ cigsd = 0.075 dlcig = 0 nigc = 1
+ poxedge = 1 pigcd = 1 ntox = 1
+ toxref = 4.23E-9 agidl = 0 bgidl = 2.3E9
+ cgidl = 0.5 egidl = 0.8 noia = 3E41
+ noib = 0 noic = 0 em = 4.1E7
+ af = 1 ef = 0.88 kf = 0
+ lintnoi = 0 tnoia = 2.5E7 tnoib = 0
+ ntnoi = 1 rnoia = 0.69 rnoib = 0.34
+ xpart = 0 cgso = {2E-11/sw_func_tox_lv_ratio} cgdo = {2E-11/sw_func_tox_lv_ratio}
+ cgbo = {1E-13/sw_func_tox_lv_ratio} ckappas = 0.6 cf = 0
+ clc = 7E-8 cle = 0.492 dlc = -1.2E-8
+ dwc = 0 vfbcv = -1 noff = 2.6123
+ voffcv = 0.112 acde = 0.44 moin = 8.7
+ cgsl = {0/sw_func_tox_lv_ratio} cgdl = {0/sw_func_tox_lv_ratio} ijthsrev = 0.1
+ ijthsfwd = 0.1 xjbvs = 1 bvs = 12.69
+ jss = 2.1483E-5 jsws = 1.4472E-10 cjs = {7.682E-04*sw_func_psd_nw_cj}
+ mjs = 0.3362 mjsws = 0.2659 cjsws = {9.160236799999998E-11*sw_func_psd_nw_cj}
+ cjswgs = {2.39155046E-10*sw_func_psd_nw_cj} mjswgs = 0.9274 pbs = 0.6587
+ pbsws = 0.7418 pbswgs = 1.4338 xrcrg1 = 12
+ xrcrg2 = 1 rbpb = 50 rbpd = 50
+ rbps = 50 rbdb = 50 rbsb = 50
+ gbmin = 1E-12 tnom = 30 ute = -0.130799664204516
+ lute = -1.855454574248183E-7 wute = 1.87553929252976E-8 pute = 9.927572590423421E-14
+ kt1 = -0.528071656533333 wkt1 = -6.233220567515299E-8 kt1l = 0
+ kt2 = -0.055045 ua1 = 6.9609E-10 ub1 = 9.658631218199466E-20
+ lub1 = -4.3570921301577E-25 wub1 = -1.168899634003519E-25 pub1 = 2.331253430056617E-31
+ uc1 = -9.961E-12 at = 3.008993546731378E5 lat = -0.102334997726826
+ wat = 2.887468569230978E-3 pat = -2.439906233454626E-8 prt = 0
+ njs = 1.3632 xtis = 5.2 tpb = 1.671E-3
+ tpbsw = 1.246E-3 tpbswg = 0 tcj = 1.2407E-3
+ tcjsw = 3.7357E-4 tcjswg = 2E-12 tvoff = 0
+ tvfbsdoff = 0 saref = 3E-6 sbref = 3E-6
+ wlod = 0 ku0 = 5.9E-8 kvsat = 0
+ kvth0 = 1.76E-8 tku0 = 0 llodku0 = 0
+ wlodku0 = 1 llodvth = 0 wlodvth = 1
+ lku0 = 0 wku0 = 0 pku0 = 0
+ lkvth0 = 0 wkvth0 = 7.3E-7 pkvth0 = 0
+ stk2 = 0 lodk2 = 1 steta0 = 0
+ lodeta0 = 1

.model plowvt_model.32 pmos
+ level = 54 lmin = 1.5E-6 lmax = 2E-6 wmin = 5.5E-7
+ wmax = 1E-6 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 4.23E-9
+ toxm = 4.23E-9 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 9.999999999999999E22 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {7.476E-9+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {2.8E-9-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = -7.916E-9 dwb = 0 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = -0.670211763626513 lvth0 = 4.585943712804615E-7
+ wvth0 = 1.911501046471693E-7 pvth0 = -2.887967969991329E-13 k1 = 0.64774
+ k2 = -0.142600147982282 lk2 = 1.623882710603925E-7 wk2 = 7.741440016406353E-8
+ pk2 = -1.16476925267449E-13 k3 = 3.39 k3b = 1
+ w0 = 1E-8 lpe0 = 0 lpeb = 0
+ vbm = -3 dvtp0 = 0 dvtp1 = 0
+ dvt0 = 2.4422 dvt1 = 0.16136 dvt2 = 0.026237
+ dvt0w = 0.5 dvt1w = 1.9281E6 dvt2w = -0.032
+ vfbsdoff = 0 u0 = 5.79942163890759E-3 lu0 = -5.136686490834932E-9
+ wu0 = -3.083330826343265E-9 pu0 = 5.063065235282099E-15 ua = -1.543688882016711E-9
+ lua = -2.216242263280271E-15 wua = -1.322536396547203E-15 pua = 2.183105008959705E-21
+ ub = 1.570149107783111E-18 lub = 2.384923318176564E-24 wub = 1.371532461676462E-24
+ pub = -2.349263944723188E-30 uc = 1.417233802938311E-10 luc = -1.303025711877448E-16
+ wuc = -7.598402218367774E-17 puc = 1.283542871433456E-22 ud = 0
+ up = 0 lp = 1 eu = 1.67
+ vsat = 1.612644557073066E4 lvsat = 0.214664360953735 wvsat = 0.106024217523443
+ pvsat = -2.114546994287545E-7 a0 = 0.312723262515484 la0 = 1.72389672717115E-6
+ wa0 = 1.329713412441775E-6 pa0 = -2.105296549334326E-12 ags = 0.706329809819307
+ lags = -4.787866901897053E-7 wags = -4.484558069711124E-7 pags = 7.373826384596227E-13
+ b0 = 4.082320739876978E-7 lb0 = -5.651169710989845E-13 wb0 = -4.021281880174337E-13
+ pb0 = 5.566673421471124E-19 b1 = 2.580668054468268E-7 lb1 = -9.959978422090713E-13
+ wb1 = -2.542081905717858E-13 pb1 = 9.811056824723614E-19 keta = -9.896979213084448E-3
+ lketa = -5.351016657424376E-9 wketa = -2.64290426010959E-9 pketa = 5.271008256362566E-15
+ a1 = 0 a2 = 0.46703705 rdsw = 484.7
+ rdswmin = 0 rdw = 0 rdwmin = 0
+ rsw = 0 rswmin = 0 prwb = 0.1
+ prwg = 0.052 wr = 1 voff = -0.1819
+ voffl = 0 minv = 0 nfactor = 2.5373
+ eta0 = 0.2 etab = -2.5E-4 dsub = 1
+ cit = -6.393105E-11 cdsc = 2.8125E-7 cdscb = 1E-4
+ cdscd = 1E-10 pclm = 0.030097 pdiblc1 = 0
+ pdiblc2 = 1.502160855295993E-3 lpdiblc2 = 2.000595258398966E-8 wpdiblc2 = -1.780428732588169E-8
+ ppdiblc2 = 3.084412513458259E-14 pdiblcb = -0.025 drout = 0.43496
+ pscbe1 = 8E8 pscbe2 = 8.6797E-9 pvag = 0
+ delta = -0.100843198228025 ldelta = 2.479227799089169E-7 wdelta = 5.619743110817708E-8
+ pdelta = -1.109215618239584E-13 fprout = 0 pdits = 0
+ pditsl = 0 pditsd = 0 lambda = 0
+ vtl = 0 lc = 5E-9 xn = 3
+ alpha0 = 5.0449517E-13 alpha1 = -4.0583656E-18 beta0 = 6.2016506
+ aigbacc = 0.43 bigbacc = 0.054 cigbacc = 0.075
+ nigbacc = 1 aigbinv = 0.35 bigbinv = 0.03
+ cigbinv = 6E-3 eigbinv = 1.1 nigbinv = 3
+ aigc = 0.43 bigc = 0.054 cigc = 0.075
+ aigsd = 0.43 bigsd = 0.054 cigsd = 0.075
+ dlcig = 0 nigc = 1 poxedge = 1
+ pigcd = 1 ntox = 1 toxref = 4.23E-9
+ agidl = 0 bgidl = 2.3E9 cgidl = 0.5
+ egidl = 0.8 noia = 3E41 noib = 0
+ noic = 0 em = 4.1E7 af = 1
+ ef = 0.88 kf = 0 lintnoi = 0
+ tnoia = 2.5E7 tnoib = 0 ntnoi = 1
+ rnoia = 0.69 rnoib = 0.34 xpart = 0
+ cgso = {2E-11/sw_func_tox_lv_ratio} cgdo = {2E-11/sw_func_tox_lv_ratio} cgbo = {1E-13/sw_func_tox_lv_ratio}
+ ckappas = 0.6 cf = 0 clc = 7E-8
+ cle = 0.492 dlc = -1.2E-8 dwc = 0
+ vfbcv = -1 noff = 2.6123 voffcv = 0.112
+ acde = 0.44 moin = 8.7 cgsl = {0/sw_func_tox_lv_ratio}
+ cgdl = {0/sw_func_tox_lv_ratio} ijthsrev = 0.1 ijthsfwd = 0.1
+ xjbvs = 1 bvs = 12.69 jss = 2.1483E-5
+ jsws = 1.4472E-10 cjs = {7.682E-04*sw_func_psd_nw_cj} mjs = 0.3362
+ mjsws = 0.2659 cjsws = {9.160236799999998E-11*sw_func_psd_nw_cj} cjswgs = {2.39155046E-10*sw_func_psd_nw_cj}
+ mjswgs = 0.9274 pbs = 0.6587 pbsws = 0.7418
+ pbswgs = 1.4338 xrcrg1 = 12 xrcrg2 = 1
+ rbpb = 50 rbpd = 50 rbps = 50
+ rbdb = 50 rbsb = 50 gbmin = 1E-12
+ tnom = 30 ute = -0.208920260845853 lute = -2.974173948333561E-8
+ wute = 6.735645223810137E-8 pute = 2.345773210778403E-15 kt1 = -0.122598227245512
+ lkt1 = -8.086762073716319E-7 wkt1 = -3.854316271428555E-7 pkt1 = 6.443894861751859E-13
+ kt1l = 0 kt2 = -0.288747101858987 lkt2 = 4.660954719475632E-7
+ wkt2 = 1.734865365973928E-7 pkt2 = -3.460015485898401E-13 ua1 = 1.14980393757184E-9
+ lua1 = -9.04887077093278E-16 wua1 = -2.860637564717299E-16 pua1 = 5.705255559072181E-22
+ ub1 = -7.484405044242205E-19 lub1 = 1.249612270023665E-24 wub1 = 2.905724461234136E-25
+ pub1 = -5.79517686548536E-31 uc1 = 1.320472035310364E-10 luc1 = -2.83221161122299E-16
+ wuc1 = -1.398848968718404E-16 puc1 = 2.789864383211985E-22 at = 3.130523743601778E5
+ lat = -0.126572980190659 wat = 0.150978206130312 pat = -3.197512293263655E-7
+ prt = 0 njs = 1.3632 xtis = 5.2
+ tpb = 1.671E-3 tpbsw = 1.246E-3 tpbswg = 0
+ tcj = 1.2407E-3 tcjsw = 3.7357E-4 tcjswg = 2E-12
+ tvoff = 0 tvfbsdoff = 0 saref = 3E-6
+ sbref = 3E-6 wlod = 0 ku0 = 5.9E-8
+ kvsat = 0 kvth0 = 1.76E-8 tku0 = 0
+ llodku0 = 0 wlodku0 = 1 llodvth = 0
+ wlodvth = 1 lku0 = 0 wku0 = 0
+ pku0 = 0 lkvth0 = 0 wkvth0 = 7.3E-7
+ pkvth0 = 0 stk2 = 0 lodk2 = 1
+ steta0 = 0 lodeta0 = 1

.model plowvt_model.33 pmos
+ level = 54 lmin = 1E-6 lmax = 1.5E-6 wmin = 5.5E-7
+ wmax = 1E-6 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 4.23E-9
+ toxm = 4.23E-9 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 9.999999999999999E22 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {7.476E-9+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {2.8E-9-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = -7.916E-9 dwb = 0 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = -0.363336515178667 wvth0 = -2.102570004284754E-9
+ k1 = 0.64774 k2 = -0.033935619703111 wk2 = -5.278678146898043E-10
+ k3 = 3.39 k3b = 1 w0 = 1E-8
+ lpe0 = 0 lpeb = 0 vbm = -3
+ dvtp0 = 0 dvtp1 = 0 dvt0 = 2.4422
+ dvt1 = 0.16136 dvt2 = 0.026237 dvt0w = 0.5
+ dvt1w = 1.9281E6 dvt2w = -0.032 vfbsdoff = 0
+ u0 = 2.362131428231111E-3 wu0 = 3.046946255318006E-10 ua = -3.026720375111111E-9
+ wua = 1.383208096624496E-16 ub = 3.166056039111111E-18 wub = -2.005124692143217E-25
+ uc = 5.452947559111111E-11 wuc = 9.906159255927181E-18 ud = 0
+ up = 0 lp = 1 eu = 1.67
+ vsat = 1.597722973866667E5 wvsat = -0.035473841516141 a0 = 1.466294412924445
+ wa0 = -7.907710504639821E-8 ags = 0.385942570666667 wags = 4.497475944994132E-8
+ b0 = 3.007564257777778E-8 wb0 = -2.962595156995484E-14 b1 = -4.084199733333335E-7
+ wb1 = 4.023132778920534E-13 keta = -0.013477691644444 wketa = 8.842693589767097E-10
+ a1 = 0 a2 = 0.46703705 rdsw = 484.7
+ rdswmin = 0 rdw = 0 rdwmin = 0
+ rsw = 0 rswmin = 0 prwb = 0.1
+ prwg = 0.052 wr = 1 voff = -0.1819
+ voffl = 0 minv = 0 nfactor = 2.5373
+ eta0 = 0.2 etab = -2.5E-4 dsub = 1
+ cit = -6.393105E-11 cdsc = 2.8125E-7 cdscb = 1E-4
+ cdscd = 1E-10 pclm = 0.030097 pdiblc1 = 0
+ pdiblc2 = 0.01488944176 wpdiblc2 = 2.83551803719552E-9 pdiblcb = -0.025
+ drout = 0.43496 pscbe1 = 8E8 pscbe2 = 8.6797E-9
+ pvag = 0 delta = 0.065058019591111 wdelta = -1.802738274618482E-8
+ fprout = 0 pdits = 0 pditsl = 0
+ pditsd = 0 lambda = 0 vtl = 0
+ lc = 5E-9 xn = 3 alpha0 = 5.0449517E-13
+ alpha1 = -4.0583656E-18 beta0 = 6.2016506 aigbacc = 0.43
+ bigbacc = 0.054 cigbacc = 0.075 nigbacc = 1
+ aigbinv = 0.35 bigbinv = 0.03 cigbinv = 6E-3
+ eigbinv = 1.1 nigbinv = 3 aigc = 0.43
+ bigc = 0.054 cigc = 0.075 aigsd = 0.43
+ bigsd = 0.054 cigsd = 0.075 dlcig = 0
+ nigc = 1 poxedge = 1 pigcd = 1
+ ntox = 1 toxref = 4.23E-9 agidl = 0
+ bgidl = 2.3E9 cgidl = 0.5 egidl = 0.8
+ noia = 3E41 noib = 0 noic = 0
+ em = 4.1E7 af = 1 ef = 0.88
+ kf = 0 lintnoi = 0 tnoia = 2.5E7
+ tnoib = 0 ntnoi = 1 rnoia = 0.69
+ rnoib = 0.34 xpart = 0 cgso = {2E-11/sw_func_tox_lv_ratio}
+ cgdo = {2E-11/sw_func_tox_lv_ratio} cgbo = {1E-13/sw_func_tox_lv_ratio} ckappas = 0.6
+ cf = 0 clc = 7E-8 cle = 0.492
+ dlc = -1.2E-8 dwc = 0 vfbcv = -1
+ noff = 2.6123 voffcv = 0.112 acde = 0.44
+ moin = 8.7 cgsl = {0/sw_func_tox_lv_ratio} cgdl = {0/sw_func_tox_lv_ratio}
+ ijthsrev = 0.1 ijthsfwd = 0.1 xjbvs = 1
+ bvs = 12.69 jss = 2.1483E-5 jsws = 1.4472E-10
+ cjs = {7.682E-04*sw_func_psd_nw_cj} mjs = 0.3362 mjsws = 0.2659
+ cjsws = {9.160236799999998E-11*sw_func_psd_nw_cj} cjswgs = {2.39155046E-10*sw_func_psd_nw_cj} mjswgs = 0.9274
+ pbs = 0.6587 pbsws = 0.7418 pbswgs = 1.4338
+ xrcrg1 = 12 xrcrg2 = 1 rbpb = 50
+ rbpd = 50 rbps = 50 rbdb = 50
+ rbsb = 50 gbmin = 1E-12 tnom = 30
+ ute = -0.228822388444444 wute = 6.89261612924231E-8 kt1 = -0.663735946311111
+ wkt1 = 4.577118748186739E-8 kt1l = 0 kt2 = 0.023147619733333
+ wkt2 = -5.804554891508053E-8 ua1 = 5.442852832E-10 wua1 = 9.571190995440641E-17
+ ub1 = 8.775614307555558E-20 wub1 = -9.722043834428986E-26 uc1 = -5.747445139555556E-11
+ wuc1 = 4.680303027028921E-17 at = 2.283541809777778E5 wat = -0.062988087583798
+ prt = 0 njs = 1.3632 xtis = 5.2
+ tpb = 1.671E-3 tpbsw = 1.246E-3 tpbswg = 0
+ tcj = 1.2407E-3 tcjsw = 3.7357E-4 tcjswg = 2E-12
+ tvoff = 0 tvfbsdoff = 0 saref = 2.74E-6
+ sbref = 2.74E-6 wlod = 0 ku0 = 5.9E-8
+ kvsat = 0 kvth0 = 1.76E-8 tku0 = 0
+ llodku0 = 0 wlodku0 = 1 llodvth = 0
+ wlodvth = 1 lku0 = 0 wku0 = 0
+ pku0 = 0 lkvth0 = 0 wkvth0 = 7.3E-7
+ pkvth0 = 0 stk2 = 0 lodk2 = 1
+ steta0 = 0 lodeta0 = 1

.model plowvt_model.34 pmos
+ level = 54 lmin = 5E-7 lmax = 1E-6 wmin = 5.5E-7
+ wmax = 1E-6 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 4.23E-9
+ toxm = 4.23E-9 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 9.999999999999999E22 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {7.476E-9+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {2.8E-9-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = -7.916E-9 dwb = 0 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = -0.401918740249668 lvth0 = 3.836616461060401E-8
+ wvth0 = 3.011322572894964E-8 pvth0 = -3.203538727712828E-14 k1 = 0.64774
+ k2 = -0.029205731136259 lk2 = -4.703401190877893E-9 wk2 = -2.832255305792256E-9
+ pk2 = 2.291482921152278E-15 k3 = 3.39 k3b = 1
+ w0 = 1E-8 lpe0 = 0 lpeb = 0
+ vbm = -3 dvtp0 = 0 dvtp1 = 0
+ dvt0 = 2.4422 dvt1 = 0.16136 dvt2 = 0.026237
+ dvt0w = 0.5 dvt1w = 1.9281E6 dvt2w = -0.032
+ vfbsdoff = 0 u0 = 2.463957687421042E-3 lu0 = -1.01256032138467E-10
+ wu0 = 2.494683081691499E-10 pu0 = 5.491704998541977E-17 ua = -3.101914626511644E-9
+ lua = 7.477316359268981E-17 wua = 2.513513751120419E-16 pua = -1.123975942830746E-22
+ ub = 3.33172836638151E-18 lub = -1.647445622376853E-25 wub = -4.416289008393744E-25
+ pub = 2.397661796079525E-31 uc = 6.494258831678579E-11 luc = -1.035479929441089E-17
+ wuc = 7.197363225326794E-18 puc = 2.693626772829024E-24 ud = 0
+ up = 0 lp = 1 eu = 1.67
+ vsat = 1.863063690625707E5 lvsat = -0.026385480874519 wvsat = -0.042922741075278
+ pvsat = 7.407185721605916E-9 a0 = 1.766488568424135 la0 = -2.985130682288924E-7
+ wa0 = -1.572685465162768E-7 pa0 = 7.775356939764723E-14 ags = 0.79921751339008
+ lags = -4.109606030441621E-7 wags = -1.920188359763355E-7 pags = 2.356664312918896E-13
+ b0 = 8.752903572209777E-8 lb0 = -5.713165414271179E-14 wb0 = 2.111620237649904E-14
+ pb0 = -5.045799788435375E-20 b1 = -5.701314861533867E-7 lb1 = 1.60805928348261E-13
+ wb1 = 4.527022113214772E-13 pb1 = -5.010675540221912E-20 keta = -0.013477691644444
+ wketa = 8.842693589767097E-10 a1 = 0 a2 = 0.46703705
+ rdsw = 484.7 rdswmin = 0 rdw = 0
+ rdwmin = 0 rsw = 0 rswmin = 0
+ prwb = 0.1 prwg = 0.052 wr = 1
+ voff = -0.1819 voffl = 0 minv = 0
+ nfactor = 2.5373 eta0 = 0.2 etab = -2.5E-4
+ dsub = 1 cit = -6.393105E-11 cdsc = 2.8125E-7
+ cdscb = 1E-4 cdscd = 1E-10 pclm = 0.030097
+ pdiblc1 = 0 pdiblc2 = 0.013003747107584 lpdiblc2 = 1.875134762362461E-9
+ wpdiblc2 = -2.625827156551621E-8 ppdiblc2 = 2.893086438093654E-14 pdiblcb = -0.025
+ drout = 0.43496 pscbe1 = 8E8 pscbe2 = 8.6797E-9
+ pvag = 0 delta = 0.036097795152156 ldelta = 2.879804718209651E-8
+ wdelta = -4.183454678721413E-9 pdelta = -1.376640207028561E-14 fprout = 0
+ pdits = 0 pditsl = 0 pditsd = 0
+ lambda = 0 vtl = 0 lc = 5E-9
+ xn = 3 alpha0 = 5.0449517E-13 alpha1 = -4.0583656E-18
+ beta0 = 6.2016506 aigbacc = 0.43 bigbacc = 0.054
+ cigbacc = 0.075 nigbacc = 1 aigbinv = 0.35
+ bigbinv = 0.03 cigbinv = 6E-3 eigbinv = 1.1
+ nigbinv = 3 aigc = 0.43 bigc = 0.054
+ cigc = 0.075 aigsd = 0.43 bigsd = 0.054
+ cigsd = 0.075 dlcig = 0 nigc = 1
+ poxedge = 1 pigcd = 1 ntox = 1
+ toxref = 4.23E-9 agidl = 0 bgidl = 2.3E9
+ cgidl = 0.5 egidl = 0.8 noia = 3E41
+ noib = 0 noic = 0 em = 4.1E7
+ af = 1 ef = 0.88 kf = 0
+ lintnoi = 0 tnoia = 2.5E7 tnoib = 0
+ ntnoi = 1 rnoia = 0.69 rnoib = 0.34
+ xpart = 0 cgso = {2E-11/sw_func_tox_lv_ratio} cgdo = {2E-11/sw_func_tox_lv_ratio}
+ cgbo = {1E-13/sw_func_tox_lv_ratio} ckappas = 0.6 cf = 0
+ clc = 7E-8 cle = 0.492 dlc = -1.2E-8
+ dwc = 0 vfbcv = -1 noff = 2.6123
+ voffcv = 0.112 acde = 0.44 moin = 8.7
+ cgsl = {0/sw_func_tox_lv_ratio} cgdl = {0/sw_func_tox_lv_ratio} ijthsrev = 0.1
+ ijthsfwd = 0.1 xjbvs = 1 bvs = 12.69
+ jss = 2.1483E-5 jsws = 1.4472E-10 cjs = {7.682E-04*sw_func_psd_nw_cj}
+ mjs = 0.3362 mjsws = 0.2659 cjsws = {9.160236799999998E-11*sw_func_psd_nw_cj}
+ cjswgs = {2.39155046E-10*sw_func_psd_nw_cj} mjswgs = 0.9274 pbs = 0.6587
+ pbsws = 0.7418 pbswgs = 1.4338 xrcrg1 = 12
+ xrcrg2 = 1 rbpb = 50 rbpd = 50
+ rbps = 50 rbdb = 50 rbsb = 50
+ gbmin = 1E-12 tnom = 30 ute = -0.064992987668764
+ lute = -1.629119561313362E-7 wute = -1.873043193380294E-8 pute = 8.716571630415918E-14
+ kt1 = -0.658233325992391 lkt1 = -5.471805644935067E-9 wkt1 = 6.081490720717695E-8
+ pkt1 = -1.495947489484784E-14 kt1l = 0 kt2 = 0.056036875180373
+ lkt2 = -3.270507561653658E-8 wkt2 = -7.56428792635084E-8 pkt2 = 1.749878529847666E-14
+ ua1 = -7.44036427946675E-12 lua1 = 5.486359838535817E-16 wua1 = 3.909116141870001E-16
+ pua1 = -2.935465858888912E-22 ub1 = 1.221374060596452E-18 lub1 = -1.127269657182779E-24
+ wub1 = -6.058788286684615E-25 pub1 = 5.058099033383562E-31 uc1 = -8.568713393579236E-11
+ luc1 = 2.805469151801148E-17 wuc1 = 6.189816963807783E-17 puc1 = -1.5010606587329E-23
+ at = 4.406018237398472E5 lat = -0.211059055962602 wat = -0.171053878094022
+ pat = 1.074606220833664E-7 prt = 0 njs = 1.3632
+ xtis = 5.2 tpb = 1.671E-3 tpbsw = 1.246E-3
+ tpbswg = 0 tcj = 1.2407E-3 tcjsw = 3.7357E-4
+ tcjswg = 2E-12 tvoff = 0 tvfbsdoff = 0
+ saref = 2.74E-6 sbref = 2.74E-6 wlod = 0
+ ku0 = 5.9E-8 kvsat = 0 kvth0 = 1.76E-8
+ tku0 = 0 llodku0 = 0 wlodku0 = 1
+ llodvth = 0 wlodvth = 1 lku0 = 0
+ wku0 = 0 pku0 = 0 lkvth0 = 0
+ wkvth0 = 7.3E-7 pkvth0 = 0 stk2 = 0
+ lodk2 = 1 steta0 = 0 lodeta0 = 1

.model plowvt_model.35 pmos
+ level = 54 lmin = 3.5E-7 lmax = 5E-7 wmin = 5.5E-7
+ wmax = 1E-6 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 4.23E-9
+ toxm = 4.23E-9 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 9.999999999999999E22 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {7.476E-9+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {2.8E-9-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = -7.916E-9 dwb = 0 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = -0.178228999854364 lvth0 = -7.222604304083425E-8
+ wvth0 = -1.34898549039522E-7 pvth0 = 4.95464341684041E-14 k1 = 0.64774
+ k2 = -0.04695523411456 lk2 = 4.071953081594203E-9 wk2 = -1.048260449569369E-8
+ pk2 = 6.073815560639547E-15 k3 = 3.39 k3b = 1
+ w0 = 1E-8 lpe0 = 0 lpeb = 0
+ vbm = -3 dvtp0 = 0 dvtp1 = 0
+ dvt0 = 2.4422 dvt1 = 0.16136 dvt2 = 0.026237
+ dvt0w = 0.5 dvt1w = 1.9281E6 dvt2w = -0.032
+ vfbsdoff = 0 u0 = 9.335311067710586E-4 lu0 = 6.553868693348846E-10
+ wu0 = 1.170785149259878E-9 pu0 = -4.005819962498363E-16 ua = -3.076683125774223E-9
+ lua = 6.229870962810906E-17 wua = 2.386014055976464E-16 pua = -1.060940093551574E-22
+ ub = 2.612994519040001E-18 lub = 1.905974518879572E-25 wub = -8.036427329211403E-26
+ pub = 6.115694774858691E-32 uc = 1.607392219192887E-11 luc = 1.380586923771837E-17
+ wuc = 4.015260322068485E-17 puc = -1.3599443880876E-23 ud = 0
+ up = 0 lp = 1 eu = 1.67
+ vsat = 1.729186447335822E5 lvsat = -0.019766589966267 wvsat = -0.063003950556246
+ pvsat = 1.733533568899619E-8 a0 = 1.1627 ags = -0.744608098476089
+ lags = 3.523067794624718E-7 wags = 9.865926522676745E-7 pags = -3.470390884959488E-13
+ b0 = 7.894683512234669E-7 lb0 = -4.041704517265887E-13 wb0 = -7.386199122618935E-13
+ pb0 = 3.251555371928675E-19 b1 = -1.841702327854934E-6 lb1 = 7.894705524855059E-13
+ wb1 = 1.711615945168527E-12 pb1 = -6.725137054162003E-19 keta = -0.017272271660089
+ lketa = 1.87604035973461E-9 wketa = 2.914551807187235E-9 pketa = -1.003771642395284E-15
+ a1 = 0 a2 = 0.46703705 rdsw = 484.7
+ rdswmin = 0 rdw = 0 rdwmin = 0
+ rsw = 0 rswmin = 0 prwb = 0.1
+ prwg = 0.052 wr = 1 voff = -0.1819
+ voffl = 0 minv = 0 nfactor = 2.5373
+ eta0 = 0.2 etab = -2.5E-4 dsub = 1
+ cit = -6.393105E-11 cdsc = 2.8125E-7 cdscb = 1E-4
+ cdscd = 1E-10 pclm = 0.030097 pdiblc1 = 0
+ pdiblc2 = -2.703778190791151E-3 lpdiblc2 = 9.640935269879149E-9 wpdiblc2 = -4.489995143338956E-8
+ ppdiblc2 = 3.814731090761312E-14 pdiblcb = -0.025 drout = 0.43496
+ pscbe1 = 8E8 pscbe2 = 8.6797E-9 pvag = 0
+ delta = 0.150990947607182 ldelta = -2.800512739166822E-8 wdelta = -6.545113965481561E-8
+ pdelta = 1.652434138189536E-14 fprout = 0 pdits = 0
+ pditsl = 0 pditsd = 0 lambda = 0
+ vtl = 0 lc = 5E-9 xn = 3
+ alpha0 = 5.0449517E-13 alpha1 = -4.0583656E-18 beta0 = 6.2016506
+ aigbacc = 0.43 bigbacc = 0.054 cigbacc = 0.075
+ nigbacc = 1 aigbinv = 0.35 bigbinv = 0.03
+ cigbinv = 6E-3 eigbinv = 1.1 nigbinv = 3
+ aigc = 0.43 bigc = 0.054 cigc = 0.075
+ aigsd = 0.43 bigsd = 0.054 cigsd = 0.075
+ dlcig = 0 nigc = 1 poxedge = 1
+ pigcd = 1 ntox = 1 toxref = 4.23E-9
+ agidl = 0 bgidl = 2.3E9 cgidl = 0.5
+ egidl = 0.8 noia = 3E41 noib = 0
+ noic = 0 em = 4.1E7 af = 1
+ ef = 0.88 kf = 0 lintnoi = 0
+ tnoia = 2.5E7 tnoib = 0 ntnoi = 1
+ rnoia = 0.69 rnoib = 0.34 xpart = 0
+ cgso = {2E-11/sw_func_tox_lv_ratio} cgdo = {2E-11/sw_func_tox_lv_ratio} cgbo = {1E-13/sw_func_tox_lv_ratio}
+ ckappas = 0.6 cf = 0 clc = 7E-8
+ cle = 0.492 dlc = -1.2E-8 dwc = 0
+ vfbcv = -1 noff = 2.6123 voffcv = 0.112
+ acde = 0.44 moin = 8.7 cgsl = {0/sw_func_tox_lv_ratio}
+ cgdl = {0/sw_func_tox_lv_ratio} ijthsrev = 0.1 ijthsfwd = 0.1
+ xjbvs = 1 bvs = 12.69 jss = 2.1483E-5
+ jsws = 1.4472E-10 cjs = {7.682E-04*sw_func_psd_nw_cj} mjs = 0.3362
+ mjsws = 0.2659 cjsws = {9.160236799999998E-11*sw_func_psd_nw_cj} cjswgs = {2.39155046E-10*sw_func_psd_nw_cj}
+ mjswgs = 0.9274 pbs = 0.6587 pbsws = 0.7418
+ pbswgs = 1.4338 xrcrg1 = 12 xrcrg2 = 1
+ rbpb = 50 rbpd = 50 rbps = 50
+ rbdb = 50 rbsb = 50 gbmin = 1E-12
+ tnom = 30 ute = -0.812740994898489 lute = 2.067746586430396E-7
+ wute = 5.193692717072468E-7 pute = -1.788707771759758E-13 kt1 = -0.792437324726044
+ lkt1 = 6.087865132898293E-8 wkt1 = 1.276072597769805E-7 pkt1 = -4.798161400535868E-14
+ kt1l = 0 kt2 = 0.162602047150933 lkt2 = -8.539089663878143E-8
+ wkt2 = -1.326603613960126E-7 pkt2 = 4.568822846478673E-14 ua1 = 1.972651465025422E-9
+ lua1 = -4.303214165547555E-16 wua1 = -6.685325588989222E-16 pua1 = 2.302426132847888E-22
+ ub1 = -2.955731024159289E-18 lub1 = 9.37891096720459E-25 wub1 = 1.375089402964459E-24
+ pub1 = -4.735807903809597E-31 uc1 = -1.642735166656285E-10 luc1 = 6.690779913964245E-17
+ wuc1 = 1.039456565449112E-16 puc1 = -3.579888411406741E-23 at = -4.433949910101329E4
+ lat = 0.02869593404992 wat = 0.187499153743863 pat = -6.980799685728378E-8
+ prt = 0 njs = 1.3632 xtis = 5.2
+ tpb = 1.671E-3 tpbsw = 1.246E-3 tpbswg = 0
+ tcj = 1.2407E-3 tcjsw = 3.7357E-4 tcjswg = 2E-12
+ tvoff = 0 tvfbsdoff = 0 saref = 1.74E-6
+ sbref = 1.74E-6 wlod = 0 ku0 = 5.9E-8
+ kvsat = 0 kvth0 = 1.76E-8 tku0 = 0
+ llodku0 = 0 wlodku0 = 1 llodvth = 0
+ wlodvth = 1 lku0 = 0 wku0 = 0
+ pku0 = 0 lkvth0 = 0 wkvth0 = 7.3E-7
+ pkvth0 = 0 stk2 = 0 lodk2 = 1
+ steta0 = 0 lodeta0 = 1

.model plowvt_model.36 pmos
+ level = 54 lmin = 8E-6 lmax = 2.02E-5 wmin = 4.2E-7
+ wmax = 5.5E-7 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 4.23E-9
+ toxm = 4.23E-9 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 9.999999999999999E22 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {7.476E-9+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {2.8E-9-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = -7.916E-9 dwb = 0 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = -0.324360811654753 lvth0 = -4.695322723701072E-7
+ wvth0 = -2.874662466974758E-8 pvth0 = 2.512223032670811E-13 k1 = 0.64774
+ k2 = -0.015145939918332 lk2 = -9.983469731964115E-8 wk2 = -7.065983044176135E-9
+ pk2 = 5.341635513147936E-14 k3 = 3.39 k3b = 1
+ w0 = 1E-8 lpe0 = 0 lpeb = 0
+ vbm = -3 dvtp0 = 0 dvtp1 = 0
+ dvt0 = 2.4422 dvt1 = 0.16136 dvt2 = 0.026237
+ dvt0w = 0.5 dvt1w = 1.9281E6 dvt2w = -0.032
+ vfbsdoff = 0 u0 = 2.136018588299321E-3 lu0 = -1.499076810303642E-9
+ wu0 = 7.351956081562465E-11 pu0 = 8.020780491993427E-16 ua = -3.3546384E-9
+ wua = 1.733760978432001E-16 ub = 3.679898369230768E-18 wub = -3.225795666601842E-25
+ uc = 6.0125E-11 ud = 0 up = 0
+ lp = 1 eu = 1.67 vsat = 1.2376E5
+ a0 = 1.691430168333539 la0 = 7.009802692698966E-6 wa0 = 1.73729184934765E-8
+ pa0 = -3.750580911123196E-12 ags = 0.614166424 wags = -1.87029465548352E-7
+ b0 = 2.194793062540307E-7 lb0 = -3.184915681691648E-12 wb0 = -1.623203508606066E-13
+ pb0 = 1.704082765657752E-18 b1 = 1.229343754146461E-7 lb1 = 8.134525327229119E-14
+ wb1 = 4.347030894314441E-14 pb1 = -4.352361507283285E-20 keta = -0.01258
+ a1 = 0 a2 = 0.46703705 rdsw = 484.7
+ rdswmin = 0 rdw = 0 rdwmin = 0
+ rsw = 0 rswmin = 0 prwb = 0.1
+ prwg = 0.052 wr = 1 voff = -0.1819
+ voffl = 0 minv = 0 nfactor = 2.5373
+ eta0 = 0.2 etab = -2.5E-4 dsub = 1
+ cit = -6.393105E-11 cdsc = 2.8125E-7 cdscb = 1E-4
+ cdscd = 1E-10 pclm = -0.452449145415385 wpclm = 2.581853500122107E-7
+ pdiblc1 = 0 pdiblc2 = 3.630289877787937E-3 lpdiblc2 = -4.524082665026862E-8
+ wpdiblc2 = -1.71074635837068E-9 ppdiblc2 = 2.420601381757292E-14 pdiblcb = -0.025
+ drout = 0.462067058461539 wdrout = -1.45035774157293E-8 pscbe1 = 8E8
+ pscbe2 = 8.6797E-9 pvag = 0 delta = 0.021899488076812
+ ldelta = -2.316264584248252E-7 wdelta = -4.45453574452227E-9 pdelta = 1.239312733272859E-13
+ fprout = 0 pdits = 0 pditsl = 0
+ pditsd = 0 lambda = 0 vtl = 0
+ lc = 5E-9 xn = 3 alpha0 = 5.0449517E-13
+ alpha1 = -4.0583656E-18 beta0 = 6.2016506 aigbacc = 0.43
+ bigbacc = 0.054 cigbacc = 0.075 nigbacc = 1
+ aigbinv = 0.35 bigbinv = 0.03 cigbinv = 6E-3
+ eigbinv = 1.1 nigbinv = 3 aigc = 0.43
+ bigc = 0.054 cigc = 0.075 aigsd = 0.43
+ bigsd = 0.054 cigsd = 0.075 dlcig = 0
+ nigc = 1 poxedge = 1 pigcd = 1
+ ntox = 1 toxref = 4.23E-9 agidl = 0
+ bgidl = 2.3E9 cgidl = 0.5 egidl = 0.8
+ noia = 3E41 noib = 0 noic = 0
+ em = 4.1E7 af = 1 ef = 0.88
+ kf = 0 lintnoi = 0 tnoia = 2.5E7
+ tnoib = 0 ntnoi = 1 rnoia = 0.69
+ rnoib = 0.34 xpart = 0 cgso = {2E-11/sw_func_tox_lv_ratio}
+ cgdo = {2E-11/sw_func_tox_lv_ratio} cgbo = {1E-13/sw_func_tox_lv_ratio} ckappas = 0.6
+ cf = 0 clc = 7E-8 cle = 0.492
+ dlc = -1.2E-8 dwc = 0 vfbcv = -1
+ noff = 2.6123 voffcv = 0.112 acde = 0.44
+ moin = 8.7 cgsl = {0/sw_func_tox_lv_ratio} cgdl = {0/sw_func_tox_lv_ratio}
+ ijthsrev = 0.1 ijthsfwd = 0.1 xjbvs = 1
+ bvs = 12.69 jss = 2.1483E-5 jsws = 1.4472E-10
+ cjs = {7.682E-04*sw_func_psd_nw_cj} mjs = 0.3362 mjsws = 0.2659
+ cjsws = {9.160236799999998E-11*sw_func_psd_nw_cj} cjswgs = {2.39155046E-10*sw_func_psd_nw_cj} mjswgs = 0.9274
+ pbs = 0.6587 pbsws = 0.7418 pbswgs = 1.4338
+ xrcrg1 = 12 xrcrg2 = 1 rbpb = 50
+ rbpd = 50 rbps = 50 rbdb = 50
+ rbsb = 50 gbmin = 1E-12 tnom = 30
+ ute = -0.624446655384615 wute = 1.811280099102277E-7 kt1 = -0.86149523076923
+ wkt1 = 1.000246718326153E-7 kt1l = 0 kt2 = -0.055045
+ ua1 = 6.8217E-10 ub1 = -1.76437096280615E-20 lub1 = -1.059148399749425E-24
+ wub1 = -7.088652469092495E-26 pub1 = 5.666952329891304E-31 uc1 = -9.961E-12
+ at = 2.233565131369846E5 lat = 0.681474009556644 wat = 0.031489440439083
+ pat = -3.646213058652632E-7 prt = 0 njs = 1.3632
+ xtis = 5.2 tpb = 1.671E-3 tpbsw = 1.246E-3
+ tpbswg = 0 tcj = 1.2407E-3 tcjsw = 3.7357E-4
+ tcjswg = 2E-12 tvoff = 0 tvfbsdoff = 0
+ saref = 3E-6 sbref = 3E-6 wlod = 0
+ ku0 = 5.9E-8 kvsat = 0 kvth0 = 1.76E-8
+ tku0 = 0 llodku0 = 0 wlodku0 = 1
+ llodvth = 0 wlodvth = 1 lku0 = 0
+ wku0 = 0 pku0 = 0 lkvth0 = 0
+ wkvth0 = 7.3E-7 pkvth0 = 0 stk2 = 0
+ lodk2 = 1 steta0 = 0 lodeta0 = 1

.model plowvt_model.37 pmos
+ level = 54 lmin = 4E-6 lmax = 8E-6 wmin = 4.2E-7
+ wmax = 5.5E-7 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 4.23E-9
+ toxm = 4.23E-9 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 9.999999999999999E22 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {7.476E-9+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {2.8E-9-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = -7.916E-9 dwb = 0 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = -0.449207251171784 lvth0 = 5.285401037048465E-7
+ wvth0 = 3.18153416583865E-8 pvth0 = -2.32934280346554E-13 k1 = 0.64774
+ k2 = -0.044631508417279 lk2 = 1.358847314883365E-7 wk2 = 7.212464641623218E-9
+ pk2 = -6.073126704787497E-14 k3 = 3.39 k3b = 1
+ w0 = 1E-8 lpe0 = 0 lpeb = 0
+ vbm = -3 dvtp0 = 0 dvtp1 = 0
+ dvt0 = 2.4422 dvt1 = 0.16136 dvt2 = 0.026237
+ dvt0w = 0.5 dvt1w = 1.9281E6 dvt2w = -0.032
+ vfbsdoff = 0 u0 = 2.686015463176286E-3 lu0 = -5.89597182682005E-9
+ wu0 = -1.642268208723454E-10 pu0 = 2.70271772296565E-15 ua = -3.406803156185847E-9
+ lua = 4.170259268521394E-16 wua = 2.228189933027654E-16 pua = -3.952662834619489E-22
+ ub = 4.024686478376613E-18 lub = -2.756374059755542E-24 wub = -5.235141620126904E-25
+ pub = 1.606351529086075E-30 uc = 1.008054692280246E-10 luc = -3.271901221493816E-16
+ wuc = -1.890968654879932E-17 puc = 1.519712353822199E-22 ud = 0
+ up = 0 lp = 1 eu = 1.67
+ vsat = 1.2376E5 a0 = 2.92039409414523 la0 = -2.815026515810014E-6
+ wa0 = -6.21748458902617E-7 pa0 = 1.358811028332133E-12 ags = 0.722916806783754
+ lags = -8.69394060126442E-7 wags = -2.310785905941459E-7 pags = 3.52146325266095E-13
+ b0 = -1.298512292640984E-7 lb0 = -3.922276485455163E-13 wb0 = 5.895649806072453E-14
+ pb0 = -6.4892875358937E-20 b1 = 2.069423729718154E-7 lb1 = -5.902482823987426E-13
+ wb1 = -4.628341615038879E-16 pb1 = 3.076955041629674E-19 keta = -0.01258
+ a1 = 0 a2 = 0.46703705 rdsw = 484.7
+ rdswmin = 0 rdw = 0 rdwmin = 0
+ rsw = 0 rswmin = 0 prwb = 0.1
+ prwg = 0.052 wr = 1 voff = -0.1819
+ voffl = 0 minv = 0 nfactor = 2.5373
+ eta0 = 0.2 etab = -2.5E-4 dsub = 1
+ cit = -6.393105E-11 cdsc = 2.8125E-7 cdscb = 1E-4
+ cdscd = 1E-10 pclm = -0.452449145415385 wpclm = 2.581853500122107E-7
+ pdiblc1 = 0 pdiblc2 = 1.563549316335504E-3 lpdiblc2 = -2.871847590579329E-8
+ wpdiblc2 = -2.017723506577783E-9 ppdiblc2 = 2.666011193119978E-14 pdiblcb = -0.025
+ drout = 0.462067058461539 wdrout = -1.45035774157293E-8 pscbe1 = 8E8
+ pscbe2 = 8.6797E-9 pvag = 0 delta = -4.113715150313852E-3
+ ldelta = -2.366650654588787E-8 wdelta = 7.070651695733926E-9 pdelta = 3.179431485490175E-14
+ fprout = 0 pdits = 0 pditsl = 0
+ pditsd = 0 lambda = 0 vtl = 0
+ lc = 5E-9 xn = 3 alpha0 = 5.0449517E-13
+ alpha1 = -4.0583656E-18 beta0 = 6.2016506 aigbacc = 0.43
+ bigbacc = 0.054 cigbacc = 0.075 nigbacc = 1
+ aigbinv = 0.35 bigbinv = 0.03 cigbinv = 6E-3
+ eigbinv = 1.1 nigbinv = 3 aigc = 0.43
+ bigc = 0.054 cigc = 0.075 aigsd = 0.43
+ bigsd = 0.054 cigsd = 0.075 dlcig = 0
+ nigc = 1 poxedge = 1 pigcd = 1
+ ntox = 1 toxref = 4.23E-9 agidl = 0
+ bgidl = 2.3E9 cgidl = 0.5 egidl = 0.8
+ noia = 3E41 noib = 0 noic = 0
+ em = 4.1E7 af = 1 ef = 0.88
+ kf = 0 lintnoi = 0 tnoia = 2.5E7
+ tnoib = 0 ntnoi = 1 rnoia = 0.69
+ rnoib = 0.34 xpart = 0 cgso = {2E-11/sw_func_tox_lv_ratio}
+ cgdo = {2E-11/sw_func_tox_lv_ratio} cgbo = {1E-13/sw_func_tox_lv_ratio} ckappas = 0.6
+ cf = 0 clc = 7E-8 cle = 0.492
+ dlc = -1.2E-8 dwc = 0 vfbcv = -1
+ noff = 2.6123 voffcv = 0.112 acde = 0.44
+ moin = 8.7 cgsl = {0/sw_func_tox_lv_ratio} cgdl = {0/sw_func_tox_lv_ratio}
+ ijthsrev = 0.1 ijthsfwd = 0.1 xjbvs = 1
+ bvs = 12.69 jss = 2.1483E-5 jsws = 1.4472E-10
+ cjs = {7.682E-04*sw_func_psd_nw_cj} mjs = 0.3362 mjsws = 0.2659
+ cjsws = {9.160236799999998E-11*sw_func_psd_nw_cj} cjswgs = {2.39155046E-10*sw_func_psd_nw_cj} mjswgs = 0.9274
+ pbs = 0.6587 pbsws = 0.7418 pbswgs = 1.4338
+ xrcrg1 = 12 xrcrg2 = 1 rbpb = 50
+ rbpd = 50 rbps = 50 rbdb = 50
+ rbsb = 50 gbmin = 1E-12 tnom = 30
+ ute = -1.152407129851692 lute = 4.220727217079599E-6 wute = 3.62002440606581E-7
+ pute = -1.445982548758927E-12 kt1 = -0.984775012492307 lkt1 = 9.85547887006964E-7
+ wkt1 = 1.4996699047864E-7 pkt1 = -3.9925887218378E-13 kt1l = 0
+ kt2 = -0.055045 ua1 = 6.68269488E-10 lua1 = 1.111262531327999E-16
+ ub1 = -1.7834045E-19 lub1 = 2.2552562148E-25 uc1 = -9.961E-12
+ at = 3.478857935447385E5 lat = -0.314062869735103 wat = -0.028220530804765
+ pat = 1.127240882465542E-7 prt = 0 njs = 1.3632
+ xtis = 5.2 tpb = 1.671E-3 tpbsw = 1.246E-3
+ tpbswg = 0 tcj = 1.2407E-3 tcjsw = 3.7357E-4
+ tcjswg = 2E-12 tvoff = 0 tvfbsdoff = 0
+ saref = 3E-6 sbref = 3E-6 wlod = 0
+ ku0 = 5.9E-8 kvsat = 0 kvth0 = 1.76E-8
+ tku0 = 0 llodku0 = 0 wlodku0 = 1
+ llodvth = 0 wlodvth = 1 lku0 = 0
+ wku0 = 0 pku0 = 0 lkvth0 = 0
+ wkvth0 = 7.3E-7 pkvth0 = 0 stk2 = 0
+ lodk2 = 1 steta0 = 0 lodeta0 = 1

.model plowvt_model.38 pmos
+ level = 54 lmin = 2E-6 lmax = 4E-6 wmin = 4.2E-7
+ wmax = 5.5E-7 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 4.23E-9
+ toxm = 4.23E-9 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 9.999999999999999E22 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {7.476E-9+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {2.8E-9-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = -7.916E-9 dwb = 0 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = -0.35661010920256 lvth0 = 1.58670079822976E-7
+ wvth0 = -1.205685124577276E-8 pvth0 = -5.769119301018027E-14 k1 = 0.64774
+ k2 = -0.015210822924633 lk2 = 1.836674535651064E-8 wk2 = -5.480733730589172E-9
+ pk2 = -1.002955546990981E-14 k3 = 3.39 k3b = 1
+ w0 = 1E-8 lpe0 = 0 lpeb = 0
+ vbm = -3 dvtp0 = 0 dvtp1 = 0
+ dvt0 = 2.4422 dvt1 = 0.16136 dvt2 = 0.026237
+ dvt0w = 0.5 dvt1w = 1.9281E6 dvt2w = -0.032
+ vfbsdoff = 0 u0 = 1.20794731155758E-3 lu0 = 8.023598005710463E-12
+ wu0 = 4.930828487685872E-10 pu0 = 7.71599785519096E-17 ua = -3.261358213415382E-9
+ lua = -1.639393525502059E-16 wua = 1.072397848274738E-16 pua = 6.64033068717558E-23
+ ub = 3.252542285292308E-18 lub = 3.278787051004044E-25 wub = -8.8115067573079E-26
+ pub = -1.328066137435086E-31 uc = 1.88932616E-11 wuc = 1.91363867994432E-17
+ ud = 0 up = 0 lp = 1
+ eu = 1.67 vsat = 1.2376E5 a0 = 2.005615614503385
+ la0 = 8.389646432713714E-7 wa0 = -1.691905321088072E-7 pa0 = -4.488863544530607E-13
+ ags = 0.343426817137231 lags = 6.464407545176302E-7 wags = -9.952968307327303E-8
+ pags = -1.733126309352797E-13 b0 = -3.687375558242463E-7 lb0 = 5.61979894266338E-13
+ wb0 = 9.494345851338728E-14 pb0 = -2.086391901910531E-19 b1 = -6.9486883810462E-9
+ lb1 = 2.641181730691277E-13 wb1 = 1.11579241853638E-13 pb1 = -1.398453642719153E-19
+ keta = -0.01258 a1 = 0 a2 = 0.46703705
+ rdsw = 484.7 rdswmin = 0 rdw = 0
+ rdwmin = 0 rsw = 0 rswmin = 0
+ prwb = 0.1 prwg = 0.052 wr = 1
+ voff = -0.1819 voffl = 0 minv = 0
+ nfactor = 2.5373 eta0 = 0.2 etab = -2.5E-4
+ dsub = 1 cit = -6.393105E-11 cdsc = 2.8125E-7
+ cdscb = 1E-4 cdscd = 1E-10 pclm = -0.452449145415385
+ wpclm = 2.581853500122107E-7 pdiblc1 = 0 pdiblc2 = -0.016918892351601
+ lpdiblc2 = 4.510778909261318E-8 wpdiblc2 = 8.519424579723214E-9 ppdiblc2 = -1.542947238472091E-14
+ pdiblcb = -0.025 drout = 0.462067058461539 wdrout = -1.45035774157293E-8
+ pscbe1 = 8E8 pscbe2 = 8.6797E-9 pvag = 0
+ delta = -0.048487668424295 ldelta = 1.53580812411704E-7 wdelta = 3.2134910982548E-8
+ pdelta = -6.832236244034835E-14 fprout = 0 pdits = 0
+ pditsl = 0 pditsd = 0 lambda = 0
+ vtl = 0 lc = 5E-9 xn = 3
+ alpha0 = 5.0449517E-13 alpha1 = -4.0583656E-18 beta0 = 6.2016506
+ aigbacc = 0.43 bigbacc = 0.054 cigbacc = 0.075
+ nigbacc = 1 aigbinv = 0.35 bigbinv = 0.03
+ cigbinv = 6E-3 eigbinv = 1.1 nigbinv = 3
+ aigc = 0.43 bigc = 0.054 cigc = 0.075
+ aigsd = 0.43 bigsd = 0.054 cigsd = 0.075
+ dlcig = 0 nigc = 1 poxedge = 1
+ pigcd = 1 ntox = 1 toxref = 4.23E-9
+ agidl = 0 bgidl = 2.3E9 cgidl = 0.5
+ egidl = 0.8 noia = 3E41 noib = 0
+ noic = 0 em = 4.1E7 af = 1
+ ef = 0.88 kf = 0 lintnoi = 0
+ tnoia = 2.5E7 tnoib = 0 ntnoi = 1
+ rnoia = 0.69 rnoib = 0.34 xpart = 0
+ cgso = {2E-11/sw_func_tox_lv_ratio} cgdo = {2E-11/sw_func_tox_lv_ratio} cgbo = {1E-13/sw_func_tox_lv_ratio}
+ ckappas = 0.6 cf = 0 clc = 7E-8
+ cle = 0.492 dlc = -1.2E-8 dwc = 0
+ vfbcv = -1 noff = 2.6123 voffcv = 0.112
+ acde = 0.44 moin = 8.7 cgsl = {0/sw_func_tox_lv_ratio}
+ cgdl = {0/sw_func_tox_lv_ratio} ijthsrev = 0.1 ijthsfwd = 0.1
+ xjbvs = 1 bvs = 12.69 jss = 2.1483E-5
+ jsws = 1.4472E-10 cjs = {7.682E-04*sw_func_psd_nw_cj} mjs = 0.3362
+ mjsws = 0.2659 cjsws = {9.160236799999998E-11*sw_func_psd_nw_cj} cjswgs = {2.39155046E-10*sw_func_psd_nw_cj}
+ mjswgs = 0.9274 pbs = 0.6587 pbsws = 0.7418
+ pbswgs = 1.4338 xrcrg1 = 12 xrcrg2 = 1
+ rbpb = 50 rbpd = 50 rbps = 50
+ rbdb = 50 rbsb = 50 gbmin = 1E-12
+ tnom = 30 ute = -0.143358123665034 lute = 1.901818667676112E-7
+ wute = 2.547477154272904E-8 pute = -1.017564274502768E-13 kt1 = -0.692773192140062
+ lkt1 = -1.808241842080455E-7 wkt1 = 2.579102154815574E-8 pkt1 = 9.674961811214634E-14
+ kt1l = 0 kt2 = -0.055045 ua1 = 6.9609E-10
+ ub1 = -1.2188E-19 uc1 = -9.961E-12 at = 3.06296008E5
+ lat = -0.1479366303552 prt = 0 njs = 1.3632
+ xtis = 5.2 tpb = 1.671E-3 tpbsw = 1.246E-3
+ tpbswg = 0 tcj = 1.2407E-3 tcjsw = 3.7357E-4
+ tcjswg = 2E-12 tvoff = 0 tvfbsdoff = 0
+ saref = 3E-6 sbref = 3E-6 wlod = 0
+ ku0 = 5.9E-8 kvsat = 0 kvth0 = 1.76E-8
+ tku0 = 0 llodku0 = 0 wlodku0 = 1
+ llodvth = 0 wlodvth = 1 lku0 = 0
+ wku0 = 0 pku0 = 0 lkvth0 = 0
+ wkvth0 = 7.3E-7 pkvth0 = 0 stk2 = 0
+ lodk2 = 1 steta0 = 0 lodeta0 = 1

.model plowvt_model.39 pmos
+ level = 54 lmin = 1.5E-6 lmax = 2E-6 wmin = 4.2E-7
+ wmax = 5.5E-7 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 4.23E-9
+ toxm = 4.23E-9 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 9.999999999999999E22 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {7.476E-9+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {2.8E-9-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = -7.916E-9 dwb = 0 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = -0.171745157381356 lvth0 = -2.100245800892321E-7
+ wvth0 = -7.555345609108921E-8 pvth0 = 6.894643569331886E-14 k1 = 0.64774
+ k2 = 0.032594687150218 lk2 = -7.697656393677113E-8 wk2 = -1.63232459839101E-8
+ pk2 = 1.159475096811342E-14 k3 = 3.39 k3b = 1
+ w0 = 1E-8 lpe0 = 0 lpeb = 0
+ vbm = -3 dvtp0 = 0 dvtp1 = 0
+ dvt0 = 2.4422 dvt1 = 0.16136 dvt2 = 0.026237
+ dvt0w = 0.5 dvt1w = 1.9281E6 dvt2w = -0.032
+ vfbsdoff = 0 u0 = -2.51080687834191E-4 lu0 = 2.917909039992658E-9
+ wu0 = 1.539783425752711E-10 pu0 = 7.53470005703859E-16 ua = -5.072500551867074E-9
+ lua = 3.448202927257846E-15 wua = 5.65547229782894E-16 pua = -8.476450613473341E-22
+ ub = 6.084930326449233E-18 lub = -5.321036004182967E-24 wub = -1.04409219980841E-24
+ pub = 1.773794178786634E-30 uc = -1.268606984450954E-10 luc = 2.906916979139382E-16
+ wuc = 6.772135197742741E-17 puc = -9.689785455097169E-23 ud = 0
+ up = 0 lp = 1 eu = 1.67
+ vsat = 4.963376884090094E5 lvsat = -0.743068941762928 wvsat = -0.150911847534692
+ pvsat = 3.009785887231905E-7 a0 = 5.457825096812307 la0 = -6.046121948245541E-6
+ wa0 = -1.423163033795071E-6 pa0 = 2.052036402910024E-12 ags = -1.699414509759999
+ lags = 4.720683496881466E-6 wags = 8.387328797311565E-7 pags = -2.044583486192434E-12
+ b0 = -1.792498903025822E-6 lb0 = 3.40152952512516E-12 wb0 = 7.753685197716959E-13
+ pb0 = -1.565678932364624E-18 b1 = 3.770729085252916E-7 lb1 = -5.017744998008723E-13
+ wb1 = -3.178821680117123E-13 pb1 = 7.166724715635393E-19 keta = -0.021867379647015
+ lketa = 1.852274996800745E-8 wketa = 3.761834551264282E-9 pketa = -7.502602829041483E-15
+ a1 = 0 a2 = 0.46703705 rdsw = 484.7
+ rdswmin = 0 rdw = 0 rdwmin = 0
+ rsw = 0 rswmin = 0 prwb = 0.1
+ prwg = 0.052 wr = 1 voff = -0.1819
+ voffl = 0 minv = 0 nfactor = 2.5373
+ eta0 = 0.2 etab = -2.5E-4 dsub = 1
+ cit = -6.393105E-11 cdsc = 2.8125E-7 cdscb = 1E-4
+ cdscd = 1E-10 pclm = -0.452449145415385 wpclm = 2.581853500122108E-7
+ pdiblc1 = 0 pdiblc2 = -0.070344346137118 lpdiblc2 = 1.516595141224468E-7
+ wpdiblc2 = 2.063704254739517E-8 ppdiblc2 = -3.959684965944586E-14 pdiblcb = -0.025
+ drout = 0.462067058461539 wdrout = -1.45035774157293E-8 pscbe1 = 8E8
+ pscbe2 = 8.6797E-9 pvag = 0 delta = 0.014767439463877
+ ldelta = 2.742482523953304E-8 wdelta = -5.659809367599631E-9 pdelta = 7.055427825986064E-15
+ fprout = 0 pdits = 0 pditsl = 0
+ pditsd = 0 lambda = 0 vtl = 0
+ lc = 5E-9 xn = 3 alpha0 = 5.0449517E-13
+ alpha1 = -4.0583656E-18 beta0 = 6.2016506 aigbacc = 0.43
+ bigbacc = 0.054 cigbacc = 0.075 nigbacc = 1
+ aigbinv = 0.35 bigbinv = 0.03 cigbinv = 6E-3
+ eigbinv = 1.1 nigbinv = 3 aigc = 0.43
+ bigc = 0.054 cigc = 0.075 aigsd = 0.43
+ bigsd = 0.054 cigsd = 0.075 dlcig = 0
+ nigc = 1 poxedge = 1 pigcd = 1
+ ntox = 1 toxref = 4.23E-9 agidl = 0
+ bgidl = 2.3E9 cgidl = 0.5 egidl = 0.8
+ noia = 3E41 noib = 0 noic = 0
+ em = 4.1E7 af = 1 ef = 0.88
+ kf = 0 lintnoi = 0 tnoia = 2.5E7
+ tnoib = 0 ntnoi = 1 rnoia = 0.69
+ rnoib = 0.34 xpart = 0 cgso = {2E-11/sw_func_tox_lv_ratio}
+ cgdo = {2E-11/sw_func_tox_lv_ratio} cgbo = {1E-13/sw_func_tox_lv_ratio} ckappas = 0.6
+ cf = 0 clc = 7E-8 cle = 0.492
+ dlc = -1.2E-8 dwc = 0 vfbcv = -1
+ noff = 2.6123 voffcv = 0.112 acde = 0.44
+ moin = 8.7 cgsl = {0/sw_func_tox_lv_ratio} cgdl = {0/sw_func_tox_lv_ratio}
+ ijthsrev = 0.1 ijthsfwd = 0.1 xjbvs = 1
+ bvs = 12.69 jss = 2.1483E-5 jsws = 1.4472E-10
+ cjs = {7.682E-04*sw_func_psd_nw_cj} mjs = 0.3362 mjsws = 0.2659
+ cjsws = {9.160236799999998E-11*sw_func_psd_nw_cj} cjswgs = {2.39155046E-10*sw_func_psd_nw_cj} mjswgs = 0.9274
+ pbs = 0.6587 pbsws = 0.7418 pbswgs = 1.4338
+ xrcrg1 = 12 xrcrg2 = 1 rbpb = 50
+ rbpd = 50 rbps = 50 rbdb = 50
+ rbsb = 50 gbmin = 1E-12 tnom = 30
+ ute = -0.24645302376448 lute = 3.957943355259466E-7 wute = 8.743828197218713E-8
+ pute = -2.25336452650788E-13 kt1 = -1.367460731522955 lkt1 = 1.164772644337196E-6
+ wkt1 = 2.806295660457818E-7 pkt1 = -4.115003750339189E-13 kt1l = 0
+ kt2 = 0.0354977072 lkt2 = -1.8057837523968E-7 ua1 = 2.110897745112616E-10
+ lua1 = 9.672844497147398E-16 wua1 = 2.161933790455066E-16 pua1 = -4.311760751683582E-22
+ ub1 = -6.252763284810831E-19 lub1 = 1.003973637522672E-24 wub1 = 2.246737001133897E-25
+ pub1 = -4.480892275061444E-31 uc1 = -1.293964368E-10 luc1 = 2.3820203515392E-16
+ at = 1.35111398679237E6 lat = -2.231721607258701 wat = -0.404434583478308
+ pat = 8.066043332891366E-7 prt = 0 njs = 1.3632
+ xtis = 5.2 tpb = 1.671E-3 tpbsw = 1.246E-3
+ tpbswg = 0 tcj = 1.2407E-3 tcjsw = 3.7357E-4
+ tcjswg = 2E-12 tvoff = 0 tvfbsdoff = 0
+ saref = 3E-6 sbref = 3E-6 wlod = 0
+ ku0 = 5.9E-8 kvsat = 0 kvth0 = 1.76E-8
+ tku0 = 0 llodku0 = 0 wlodku0 = 1
+ llodvth = 0 wlodvth = 1 lku0 = 0
+ wku0 = 0 pku0 = 0 lkvth0 = 0
+ wkvth0 = 7.3E-7 pkvth0 = 0 stk2 = 0
+ lodk2 = 1 steta0 = 0 lodeta0 = 1

.model plowvt_model.40 pmos
+ level = 54 lmin = 1E-6 lmax = 1.5E-6 wmin = 4.2E-7
+ wmax = 5.5E-7 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 4.23E-9
+ toxm = 4.23E-9 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 9.999999999999999E22 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {7.476E-9+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {2.8E-9-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = -7.916E-9 dwb = 0 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = -0.312286230781538 wvth0 = -2.941692257039939E-8
+ k1 = 0.64774 k2 = -0.018915326190769 wk2 = -8.564445817881305E-9
+ k3 = 3.39 k3b = 1 w0 = 1E-8
+ lpe0 = 0 lpeb = 0 vbm = -3
+ dvtp0 = 0 dvtp1 = 0 dvt0 = 2.4422
+ dvt1 = 0.16136 dvt2 = 0.026237 dvt0w = 0.5
+ dvt1w = 1.9281E6 dvt2w = -0.032 vfbsdoff = 0
+ u0 = 1.701481571261538E-3 wu0 = 6.581740102036564E-10 ua = -2.7692E-9
+ ub = 2.524279895384615E-18 wub = 1.428685729342527E-25 uc = 6.765997735384615E-11
+ wuc = 2.880710548779321E-18 ud = 0 up = 0
+ lp = 1 eu = 1.67 vsat = -897.9524923076824
+ wvsat = 0.050492454341104 a0 = 1.411972615384616 wa0 = -5.001233591630774E-8
+ ags = 1.459501106461538 wags = -5.294305880100332E-7 b0 = 4.836852010461539E-7
+ wb0 = -2.723288386093425E-13 b1 = 4.130303446153859E-8 wb1 = 1.616898820174227E-13
+ keta = -9.47260584615385E-3 wketa = -1.258643787227075E-9 a1 = 0
+ a2 = 0.46703705 rdsw = 484.7 rdswmin = 0
+ rdw = 0 rdwmin = 0 rsw = 0
+ rswmin = 0 prwb = 0.1 prwg = 0.052
+ wr = 1 voff = -0.1819 voffl = 0
+ minv = 0 nfactor = 2.5373 eta0 = 0.2
+ etab = -2.5E-4 dsub = 1 cit = -6.393105E-11
+ cdsc = 2.8125E-7 cdscb = 1E-4 cdscd = 1E-10
+ pclm = -0.452449145415385 wpclm = 2.581853500122108E-7 pdiblc1 = 0
+ pdiblc2 = 0.031140874769231 wpdiblc2 = -5.85977869152738E-9 pdiblcb = -0.025
+ drout = 0.462067058461539 wdrout = -1.45035774157293E-8 pscbe1 = 8E8
+ pscbe2 = 8.6797E-9 pvag = 0 delta = 0.033119169415385
+ wdelta = -9.385648373627035E-10 fprout = 0 pdits = 0
+ pditsl = 0 pditsd = 0 lambda = 0
+ vtl = 0 lc = 5E-9 xn = 3
+ alpha0 = 5.0449517E-13 alpha1 = -4.0583656E-18 beta0 = 6.2016506
+ aigbacc = 0.43 bigbacc = 0.054 cigbacc = 0.075
+ nigbacc = 1 aigbinv = 0.35 bigbinv = 0.03
+ cigbinv = 6E-3 eigbinv = 1.1 nigbinv = 3
+ aigc = 0.43 bigc = 0.054 cigc = 0.075
+ aigsd = 0.43 bigsd = 0.054 cigsd = 0.075
+ dlcig = 0 nigc = 1 poxedge = 1
+ pigcd = 1 ntox = 1 toxref = 4.23E-9
+ agidl = 0 bgidl = 2.3E9 cgidl = 0.5
+ egidl = 0.8 noia = 3E41 noib = 0
+ noic = 0 em = 4.1E7 af = 1
+ ef = 0.88 kf = 0 lintnoi = 0
+ tnoia = 2.5E7 tnoib = 0 ntnoi = 1
+ rnoia = 0.69 rnoib = 0.34 xpart = 0
+ cgso = {2E-11/sw_func_tox_lv_ratio} cgdo = {2E-11/sw_func_tox_lv_ratio} cgbo = {1E-13/sw_func_tox_lv_ratio}
+ ckappas = 0.6 cf = 0 clc = 7E-8
+ cle = 0.492 dlc = -1.2E-8 dwc = 0
+ vfbcv = -1 noff = 2.6123 voffcv = 0.112
+ acde = 0.44 moin = 8.7 cgsl = {0/sw_func_tox_lv_ratio}
+ cgdl = {0/sw_func_tox_lv_ratio} ijthsrev = 0.1 ijthsfwd = 0.1
+ xjbvs = 1 bvs = 12.69 jss = 2.1483E-5
+ jsws = 1.4472E-10 cjs = {7.682E-04*sw_func_psd_nw_cj} mjs = 0.3362
+ mjsws = 0.2659 cjsws = {9.160236799999998E-11*sw_func_psd_nw_cj} cjswgs = {2.39155046E-10*sw_func_psd_nw_cj}
+ mjswgs = 0.9274 pbs = 0.6587 pbsws = 0.7418
+ pbswgs = 1.4338 xrcrg1 = 12 xrcrg2 = 1
+ rbpb = 50 rbpd = 50 rbps = 50
+ rbdb = 50 rbsb = 50 gbmin = 1E-12
+ tnom = 30 ute = 0.018398646153846 wute = -6.334895882732309E-8
+ kt1 = -0.588035782153846 wkt1 = 5.267966049850978E-9 kt1l = 0
+ kt2 = -0.085339 ua1 = 8.583625593846154E-10 wua1 = -7.233450851361968E-17
+ ub1 = 4.654757243076917E-20 wub1 = -7.517187503793819E-26 uc1 = 3E-11
+ at = -1.422757396923077E5 wat = 0.13531671021089 prt = 0
+ njs = 1.3632 xtis = 5.2 tpb = 1.671E-3
+ tpbsw = 1.246E-3 tpbswg = 0 tcj = 1.2407E-3
+ tcjsw = 3.7357E-4 tcjswg = 2E-12 tvoff = 0
+ tvfbsdoff = 0 saref = 2.74E-6 sbref = 2.74E-6
+ wlod = 0 ku0 = 5.9E-8 kvsat = 0
+ kvth0 = 1.76E-8 tku0 = 0 llodku0 = 0
+ wlodku0 = 1 llodvth = 0 wlodvth = 1
+ lku0 = 0 wku0 = 0 pku0 = 0
+ lkvth0 = 0 wkvth0 = 7.3E-7 pkvth0 = 0
+ stk2 = 0 lodk2 = 1 steta0 = 0
+ lodeta0 = 1

.model plowvt_model.41 pmos
+ level = 54 lmin = 5E-7 lmax = 1E-6 wmin = 4.2E-7
+ wmax = 5.5E-7 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 4.23E-9
+ toxm = 4.23E-9 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 9.999999999999999E22 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {7.476E-9+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {2.8E-9-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = -7.916E-9 dwb = 0 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = -0.162974979299899 lvth0 = -1.484751084733421E-7
+ wvth0 = -9.773315567970242E-8 pvth0 = 6.793366220389092E-14 k1 = 0.64774
+ k2 = 0.018195764748032 lk2 = -3.690326882954394E-8 wk2 = -2.819433087569031E-8
+ pk2 = 1.951995770148527E-14 k3 = 3.39 k3b = 1
+ w0 = 1E-8 lpe0 = 0 lpeb = 0
+ vbm = -3 dvtp0 = 0 dvtp1 = 0
+ dvt0 = 2.4422 dvt1 = 0.16136 dvt2 = 0.026237
+ dvt0w = 0.5 dvt1w = 1.9281E6 dvt2w = -0.032
+ vfbsdoff = 0 u0 = 5.449906252407155E-4 lu0 = 1.150014596723106E-9
+ wu0 = 1.276207796854609E-9 pu0 = -6.145727974457074E-16 ua = -2.759653720044308E-9
+ lua = -5.400115163324527E-18 wua = 6.822536162850723E-17 pua = -6.950104183122662E-23
+ ub = 2.124083668509537E-18 lub = 3.979551280045774E-25 wub = 2.045189794676293E-25
+ pub = -6.13051642567897E-32 uc = 8.818359686399999E-11 luc = -2.040868724089697E-17
+ wuc = -5.237691915843072E-18 puc = 8.072939410820507E-24 ud = 0
+ up = 0 lp = 1 eu = 1.67
+ vsat = 1.353921310968123E5 lvsat = -0.135526859121021 wvsat = -0.015681179880175
+ pvsat = 6.580306186964032E-8 a0 = 3.281140971677539 la0 = -1.858701013497682E-6
+ wa0 = -9.676802855722036E-7 pa0 = 9.125290091378228E-13 ags = 1.337411384369231
+ lags = 1.214060196485909E-7 wags = -4.799783902559881E-7 pags = -4.917526544662244E-14
+ b0 = 1.107522024588899E-6 lb0 = -6.203433373309051E-13 wb0 = -5.24629006330705E-13
+ pb0 = 2.508872867821228E-19 b1 = -9.415855485666457E-7 lb1 = 9.773844069632267E-13
+ wb1 = 6.514479645075668E-13 pb1 = -4.870154372281992E-19 keta = -9.47260584615385E-3
+ wketa = -1.258643787227075E-9 a1 = 0 a2 = 0.46703705
+ rdsw = 484.7 rdswmin = 0 rdw = 0
+ rdwmin = 0 rsw = 0 rswmin = 0
+ prwb = 0.1 prwg = 0.052 wr = 1
+ voff = -0.1819 voffl = 0 minv = 0
+ nfactor = 2.5373 eta0 = 0.2 etab = -2.5E-4
+ dsub = 1 cit = -6.393105E-11 cdsc = 2.8125E-7
+ cdscb = 1E-4 cdscd = 1E-10 pclm = -0.828560217183015
+ lpclm = 3.740048497657321E-7 wpclm = 4.59422826739338E-7 ppclm = -2.001105468574554E-13
+ pdiblc1 = 0 pdiblc2 = -0.125264126317785 lpdiblc2 = 1.555291330809281E-7
+ wpdiblc2 = 4.772167757498043E-8 ppdiblc2 = -5.328140011141537E-14 pdiblcb = -0.025
+ drout = 0.462067058461539 wdrout = -1.45035774157293E-8 pscbe1 = 8E8
+ pscbe2 = 8.6797E-9 pvag = 0 delta = 0.094241273752911
+ ldelta = -6.077982055323598E-8 wdelta = -3.529300661709779E-8 pdelta = 3.416205690576857E-14
+ fprout = 0 pdits = 0 pditsl = 0
+ pditsd = 0 lambda = 0 vtl = 0
+ lc = 5E-9 xn = 3 alpha0 = 5.0449517E-13
+ alpha1 = -4.0583656E-18 beta0 = 6.2016506 aigbacc = 0.43
+ bigbacc = 0.054 cigbacc = 0.075 nigbacc = 1
+ aigbinv = 0.35 bigbinv = 0.03 cigbinv = 6E-3
+ eigbinv = 1.1 nigbinv = 3 aigc = 0.43
+ bigc = 0.054 cigc = 0.075 aigsd = 0.43
+ bigsd = 0.054 cigsd = 0.075 dlcig = 0
+ nigc = 1 poxedge = 1 pigcd = 1
+ ntox = 1 toxref = 4.23E-9 agidl = 0
+ bgidl = 2.3E9 cgidl = 0.5 egidl = 0.8
+ noia = 3E41 noib = 0 noic = 0
+ em = 4.1E7 af = 1 ef = 0.88
+ kf = 0 lintnoi = 0 tnoia = 2.5E7
+ tnoib = 0 ntnoi = 1 rnoia = 0.69
+ rnoib = 0.34 xpart = 0 cgso = {2E-11/sw_func_tox_lv_ratio}
+ cgdo = {2E-11/sw_func_tox_lv_ratio} cgbo = {1E-13/sw_func_tox_lv_ratio} ckappas = 0.6
+ cf = 0 clc = 7E-8 cle = 0.492
+ dlc = -1.2E-8 dwc = 0 vfbcv = -1
+ noff = 2.6123 voffcv = 0.112 acde = 0.44
+ moin = 8.7 cgsl = {0/sw_func_tox_lv_ratio} cgdl = {0/sw_func_tox_lv_ratio}
+ ijthsrev = 0.1 ijthsfwd = 0.1 xjbvs = 1
+ bvs = 12.69 jss = 2.1483E-5 jsws = 1.4472E-10
+ cjs = {7.682E-04*sw_func_psd_nw_cj} mjs = 0.3362 mjsws = 0.2659
+ cjsws = {9.160236799999998E-11*sw_func_psd_nw_cj} cjswgs = {2.39155046E-10*sw_func_psd_nw_cj} mjswgs = 0.9274
+ pbs = 0.6587 pbsws = 0.7418 pbswgs = 1.4338
+ xrcrg1 = 12 xrcrg2 = 1 rbpb = 50
+ rbpd = 50 rbps = 50 rbdb = 50
+ rbsb = 50 gbmin = 1E-12 tnom = 30
+ ute = 0.135471227470769 lute = -1.164169748615483E-7 wute = -1.259884093157802E-7
+ pute = 6.22886695657217E-14 kt1 = -0.459772642731323 lkt1 = -1.275448658417572E-7
+ wkt1 = -4.537108445029128E-8 pkt1 = 5.035547181734146E-14 kt1l = 0
+ kt2 = -0.085339 ua1 = 9.029117574331076E-10 lua1 = -4.429972253942065E-17
+ wua1 = -9.617046783106934E-17 pua1 = 2.370247794527194E-23 ub1 = 8.905531727237907E-19
+ lub1 = -8.392791689313807E-25 wub1 = -4.288737742539699E-25 pub1 = 3.51721168580422E-31
+ uc1 = 3E-11 at = -3.012027962692922E5 lat = 0.158037065060153
+ wat = 0.225847200232628 pat = -9.002351927761673E-8 prt = 0
+ njs = 1.3632 xtis = 5.2 tpb = 1.671E-3
+ tpbsw = 1.246E-3 tpbswg = 0 tcj = 1.2407E-3
+ tcjsw = 3.7357E-4 tcjswg = 2E-12 tvoff = 0
+ tvfbsdoff = 0 saref = 2.74E-6 sbref = 2.74E-6
+ wlod = 0 ku0 = 5.9E-8 kvsat = 0
+ kvth0 = 1.76E-8 tku0 = 0 llodku0 = 0
+ wlodku0 = 1 llodvth = 0 wlodvth = 1
+ lku0 = 0 wku0 = 0 pku0 = 0
+ lkvth0 = 0 wkvth0 = 7.3E-7 pkvth0 = 0
+ stk2 = 0 lodk2 = 1 steta0 = 0
+ lodeta0 = 1

.model plowvt_model.42 pmos
+ level = 54 lmin = 3.5E-7 lmax = 5E-7 wmin = 4.2E-7
+ wmax = 5.5E-7 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 4.23E-9
+ toxm = 4.23E-9 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 9.999999999999999E22 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {7.476E-9+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {2.8E-9-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = -7.916E-9 dwb = 0 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = -0.312036859599753 lvth0 = -7.477891485309417E-8
+ wvth0 = -6.330492129847108E-8 pvth0 = 5.091234312581015E-14 k1 = 0.64774
+ k2 = -0.035849167323372 lk2 = -1.018345441344165E-8 wk2 = -1.642488332018509E-8
+ pk2 = 1.370114283004349E-14 k3 = 3.39 k3b = 1
+ w0 = 1E-8 lpe0 = 0 lpeb = 0
+ vbm = -3 dvtp0 = 0 dvtp1 = 0
+ dvt0 = 2.4422 dvt1 = 0.16136 dvt2 = 0.026237
+ dvt0w = 0.5 dvt1w = 1.9281E6 dvt2w = -0.032
+ vfbsdoff = 0 u0 = 2.842284074724426E-3 lu0 = 1.423271529836022E-11
+ wu0 = 1.495106912623652E-10 pu0 = -5.7533748440902E-17 ua = -2.073443004061539E-9
+ lua = -3.446626931452058E-16 wua = -2.981802150444818E-16 pua = 1.116498752758991E-22
+ ub = 1.320790852086156E-18 lub = 7.951030964442969E-25 wub = 6.110267143042067E-25
+ pub = -2.622825883599935E-31 uc = 7.979688230400001E-11 luc = -1.626229556243298E-17
+ wuc = 6.057760858641412E-18 puc = 2.488467559115378E-24 ud = 0
+ up = 0 lp = 1 eu = 1.67
+ vsat = -4.914187452125538E5 lvsat = 0.17436843812633 wvsat = 0.292448441259654
+ pvsat = -8.653622282189151E-8 a0 = -0.478367550769231 wa0 = 8.780499109039753E-7
+ ags = 4.049647401801847 lags = -1.219523467370094E-6 wags = -1.578564164645034E-6
+ pags = 4.939655414113219E-13 b0 = -4.852296558276925E-7 lb0 = 1.671130934670573E-13
+ wb0 = -5.659529298518478E-14 pb0 = 1.949141890409764E-20 b1 = 3.412430078345847E-6
+ lb1 = -1.17524091898231E-12 wb1 = -1.099597090504388E-12 pb1 = 3.787012379697114E-19
+ keta = -9.47260584615385E-3 wketa = -1.258643787227075E-9 a1 = 0
+ a2 = 0.46703705 rdsw = 484.7 rdswmin = 0
+ rdw = 0 rdwmin = 0 rsw = 0
+ rswmin = 0 prwb = 0.1 prwg = 0.052
+ wr = 1 voff = -0.1819 voffl = 0
+ minv = 0 nfactor = 2.5373 eta0 = 0.2
+ etab = -2.5E-4 dsub = 1 cit = -6.393105E-11
+ cdsc = 2.8125E-7 cdscb = 1E-4 cdscd = 1E-10
+ pclm = -0.072077915876923 wpclm = 5.466848439011594E-8 pdiblc1 = 0
+ pdiblc2 = -0.075660718341908 lpdiblc2 = 1.310052081776545E-7 wpdiblc2 = -5.864486519414989E-9
+ ppdiblc2 = -2.678840058314627E-14 pdiblcb = -0.025 drout = 0.462067058461539
+ wdrout = -1.45035774157293E-8 pscbe1 = 8E8 pscbe2 = 8.6797E-9
+ pvag = 0 delta = 0.127550765678769 ldelta = -7.724803336138042E-8
+ wdelta = -5.290951719438213E-8 pdelta = 4.287165973517794E-14 fprout = 0
+ pdits = 0 pditsl = 0 pditsd = 0
+ lambda = 0 vtl = 0 lc = 5E-9
+ xn = 3 alpha0 = 5.0449517E-13 alpha1 = -4.0583656E-18
+ beta0 = 6.2016506 aigbacc = 0.43 bigbacc = 0.054
+ cigbacc = 0.075 nigbacc = 1 aigbinv = 0.35
+ bigbinv = 0.03 cigbinv = 6E-3 eigbinv = 1.1
+ nigbinv = 3 aigc = 0.43 bigc = 0.054
+ cigc = 0.075 aigsd = 0.43 bigsd = 0.054
+ cigsd = 0.075 dlcig = 0 nigc = 1
+ poxedge = 1 pigcd = 1 ntox = 1
+ toxref = 4.23E-9 agidl = 0 bgidl = 2.3E9
+ cgidl = 0.5 egidl = 0.8 noia = 3E41
+ noib = 0 noic = 0 em = 4.1E7
+ af = 1 ef = 0.88 kf = 0
+ lintnoi = 0 tnoia = 2.5E7 tnoib = 0
+ ntnoi = 1 rnoia = 0.69 rnoib = 0.34
+ xpart = 0 cgso = {2E-11/sw_func_tox_lv_ratio} cgdo = {2E-11/sw_func_tox_lv_ratio}
+ cgbo = {1E-13/sw_func_tox_lv_ratio} ckappas = 0.6 cf = 0
+ clc = 7E-8 cle = 0.492 dlc = -1.2E-8
+ dwc = 0 vfbcv = -1 noff = 2.6123
+ voffcv = 0.112 acde = 0.44 moin = 8.7
+ cgsl = {0/sw_func_tox_lv_ratio} cgdl = {0/sw_func_tox_lv_ratio} ijthsrev = 0.1
+ ijthsfwd = 0.1 xjbvs = 1 bvs = 12.69
+ jss = 2.1483E-5 jsws = 1.4472E-10 cjs = {7.682E-04*sw_func_psd_nw_cj}
+ mjs = 0.3362 mjsws = 0.2659 cjsws = {9.160236799999998E-11*sw_func_psd_nw_cj}
+ cjswgs = {2.39155046E-10*sw_func_psd_nw_cj} mjswgs = 0.9274 pbs = 0.6587
+ pbsws = 0.7418 pbswgs = 1.4338 xrcrg1 = 12
+ xrcrg2 = 1 rbpb = 50 rbpd = 50
+ rbps = 50 rbdb = 50 rbsb = 50
+ gbmin = 1E-12 tnom = 30 ute = 0.1579556
+ lute = -1.2753324864E-7 kt1 = -0.901871976054154 lkt1 = 9.102904455305067E-8
+ wkt1 = 1.86160051100783E-7 pkt1 = -6.411352159910967E-14 kt1l = 0
+ kt2 = -0.085339 ua1 = 1.020267348903385E-9 lua1 = -1.023203269623257E-16
+ wua1 = -1.589613423360583E-16 pua1 = 5.474628630053846E-23 ub1 = -2.126180082244924E-18
+ lub1 = 6.521937523251516E-25 wub1 = 9.312398305950617E-25 pub1 = -3.207189976569392E-31
+ uc1 = 3E-11 at = 3.651974523076924E4 lat = -8.932959457476915E-3
+ wat = 0.144235576782631 pat = -4.967473264393825E-8 prt = 0
+ njs = 1.3632 xtis = 5.2 tpb = 1.671E-3
+ tpbsw = 1.246E-3 tpbswg = 0 tcj = 1.2407E-3
+ tcjsw = 3.7357E-4 tcjswg = 2E-12 tvoff = 0
+ tvfbsdoff = 0 saref = 1.74E-6 sbref = 1.74E-6
+ wlod = 0 ku0 = 5.9E-8 kvsat = 0
+ kvth0 = 1.76E-8 tku0 = 0 llodku0 = 0
+ wlodku0 = 1 llodvth = 0 wlodvth = 1
+ lku0 = 0 wku0 = 0 pku0 = 0
+ lkvth0 = 0 wkvth0 = 7.3E-7 pkvth0 = 0
+ stk2 = 0 lodk2 = 1 steta0 = 0
+ lodeta0 = 1

.ends sky130_fd_pr__pfet_01v8_lvt
