* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

******************************************************************
******************************************************************
*  *****************************************************
*  04/24/2021 Usman Suriono
*      Why     : New scalable sky130_fd_pr__pfet_01v8 high VT model
*      What    : Converted from discrete phighvt models
*                Replaced rsh from 1 to calculated rsh from the original model.
*                PDK netlist nrd/nrs = ratio of distance the middle of the contact to Gate.
*
*  *****************************************************
*
*  Pmos High VT Model
*  -----------------------------------------------------

.subckt  sky130_fd_pr__pfet_01v8_hvt  d g s b  mult=1
+ 
.param  l = 1 w = 1 nf = 1 ad = 0 as = 0 pd = 0 ps = 0 nrd = {0.14/w} nrs = {0.14/w} sa = 0 sb = 0 sd = 0
+ swx_nrds = {361*nf/w+1489}

Msky130_fd_pr__pfet_01v8_hvt  d g s b phighvt_model l = {l} w = {w} ad = {ad} as = {as} pd = {pd} ps = {ps} nrd = {nrd} nrs = {nrs} sa = {sa} sb = {sb} sd = {sd} nf = {nf}
* + deltox = 0.3*(sw_tox_lv_corner - sw_tox_lv_nom) + sw_tox_lv_mc + sw_mm_tox_lv * mismatch_factor*MC_MM_SWITCH*AGAUSS(0,1.0,1)/sqrt(l*w*mult)
* + mulu0  = sw_u0_sky130_fd_pr__pfet_01v8_hvt
+ delvto = {(sw_vth0_sky130_fd_pr__pfet_01v8_hvt+sw_vth0_sky130_fd_pr__pfet_01v8_hvt_mc)*(0.023*8/l+0.977)*(0.024*7/w+0.976)*(0.00055*56/(w*l)+0.99945)-0.0025/l+4e-4/(l*w)+sw_mm_vth0_sky130_fd_pr__pfet_01v8_hvt*mismatch_factor*MC_MM_SWITCH*AGAUSS(0,1.0,1)/sqrt(l*w*mult)}
* + mulvsat = sw_vsat_sky130_fd_pr__pfet_01v8_hvt




.model phighvt_model.1 pmos
+ level = 54 lmin = 8E-6 lmax = 2.02E-5 wmin = 7E-6
+ wmax = 1.01E-3 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 4.23E-9
+ toxm = 4.23E-9 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 9.999999999999999E22 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {9.364E-9+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {-1.176E-8-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = -5.722E-9 dwb = -1.7864E-8 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = -1.1148095 k1 = 0.43657182
+ k2 = 0.029941288 k3 = -13.778 k3b = 2
+ w0 = 0 lpe0 = 0 lpeb = 0
+ vbm = -3 dvtp0 = 0 dvtp1 = 0
+ dvt0 = 4.05 dvt1 = 0.3 dvt2 = 0.03
+ dvt0w = -4.254 dvt1w = 1.1472E6 dvt2w = -8.96E-3
+ vfbsdoff = 0 u0 = 0.012121798 ua = -2.3807897E-10
+ ub = 8.232617299999999E-19 uc = -7.7670696E-11 ud = 0
+ up = 0 lp = 1 eu = 1.67
+ vsat = 2E5 a0 = 1.4973894 ags = 0.3864062
+ b0 = 0 b1 = 0 keta = -0.013169082
+ a1 = 0 a2 = 1 rdsw = 531.92
+ rdswmin = 0 rdw = 0 rdwmin = 0
+ rsw = 0 rswmin = 0 prwb = -0.32348
+ prwg = 0.02 wr = 1 voff = -0.19592208
+ voffl = 0 minv = 0 nfactor = 2.4926776
+ eta0 = 0.08 etab = -0.07 dsub = 0.56
+ cit = 1E-5 cdsc = 0 cdscb = 0
+ cdscd = 0 pclm = 0.075489662 pdiblc1 = 0.39
+ pdiblc2 = 3.6275994E-3 pdiblcb = -9.5744039E-5 drout = 0.56
+ pscbe1 = 7.4647513E8 pscbe2 = 9.5049925E-9 pvag = 0
+ delta = 0.01 fprout = 0 pdits = 0
+ pditsl = 0 pditsd = 0 lambda = 0
+ vtl = 0 lc = 5E-9 xn = 3
+ alpha0 = 1E-10 alpha1 = 1E-10 beta0 = 4.7923891
+ aigbacc = 0.43 bigbacc = 0.054 cigbacc = 0.075
+ nigbacc = 1 aigbinv = 0.35 bigbinv = 0.03
+ cigbinv = 6E-3 eigbinv = 1.1 nigbinv = 3
+ aigc = 0.43 bigc = 0.054 cigc = 0.075
+ aigsd = 0.43 bigsd = 0.054 cigsd = 0.075
+ dlcig = 0 nigc = 1 poxedge = 1
+ pigcd = 1 ntox = 1 toxref = 4.23E-9
+ agidl = 1E-10 bgidl = 1.1544446E9 cgidl = 300
+ egidl = 0.1 noia = 1.2E41 noib = 2E25
+ noic = 0 em = 4.1E7 af = 1
+ ef = 0.88 kf = 0 lintnoi = -6E-8
+ tnoia = 1.5 tnoib = 3.5 ntnoi = 1
+ rnoia = 0.577 rnoib = 0.37 xpart = 0
+ cgso = {5.932020000000001E-11/sw_func_tox_lv_ratio} cgdo = {5.932020000000001E-11/sw_func_tox_lv_ratio} cgbo = {0/sw_func_tox_lv_ratio}
+ ckappas = 0.6 cf = 1.2E-11 clc = 1E-7
+ cle = 0.6 dlc = -2.56E-9 dwc = 0
+ vfbcv = -0.1446893 noff = 4 voffcv = -0.1375
+ acde = 0.552 moin = 14.504 cgsl = {7.513892E-12/sw_func_tox_lv_ratio}
+ cgdl = {7.513892E-12/sw_func_tox_lv_ratio} ijthsrev = 0.1 ijthsfwd = 0.1
+ xjbvs = 1 bvs = 12.8 jss = 2.17E-5
+ jsws = 8.200000000000001E-10 cjs = {7.433E-04*sw_func_psd_nw_cj} mjs = 0.34629
+ mjsws = 0.26859 cjsws = {9.2435E-11*sw_func_psd_nw_cj} cjswgs = {2.4701E-10*sw_func_psd_nw_cj}
+ mjswgs = 0.70393 pbs = 0.6587 pbsws = 0.7418
+ pbswgs = 1.3925 xrcrg1 = 12 xrcrg2 = 1
+ rbpb = 50 rbpd = 50 rbps = 50
+ rbdb = 50 rbsb = 50 gbmin = 1E-12
+ tnom = 30 ute = -0.30066 kt1 = -0.44169
+ kt1l = 0 kt2 = -0.037961 ua1 = 2.2116E-9
+ ub1 = -7.9359E-19 uc1 = 1.1985E-10 at = 0
+ prt = 0 njs = 1.2556 xtis = 2
+ tpb = 1.9551E-3 tpbsw = 1.4242E-4 tpbswg = 0
+ tcj = 1.2407E-3 tcjsw = 0 tcjswg = 2E-12
+ tvoff = 0 tvfbsdoff = 0 saref = 3E-6
+ sbref = 3E-6 wlod = 0 ku0 = 4.5E-8
+ kvsat = 0.4 kvth0 = 2.65E-8 tku0 = 0
+ llodku0 = 0 wlodku0 = 1 llodvth = 0
+ wlodvth = 1 lku0 = 0 wku0 = 2.5E-7
+ pku0 = 0 lkvth0 = 0 wkvth0 = 2.5E-7
+ pkvth0 = 0 stk2 = 0 lodk2 = 1
+ steta0 = 0 lodeta0 = 1

.model phighvt_model.2 pmos
+ level = 54 lmin = 4E-6 lmax = 8E-6 wmin = 7E-6
+ wmax = 1.01E-3 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 4.23E-9
+ toxm = 4.23E-9 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 9.999999999999999E22 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {9.364E-9+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {-1.176E-8-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = -5.722E-9 dwb = -1.7864E-8 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = -1.123204675068 lvth0 = 6.735885506159955E-8
+ k1 = 0.443495442922 lk1 = -5.555182698712548E-8 k2 = 0.02544290814608
+ lk2 = 3.609284072552418E-8 k3 = -13.778 k3b = 2
+ w0 = 0 lpe0 = 0 lpeb = 0
+ vbm = -3 dvtp0 = 0 dvtp1 = 0
+ dvt0 = 4.05 dvt1 = 0.3 dvt2 = 0.03
+ dvt0w = -4.254 dvt1w = 1.1472E6 dvt2w = -8.96E-3
+ vfbsdoff = 0 u0 = 0.01191725833728 lu0 = 1.641128074627184E-9
+ ua = -2.594257754776E-10 lua = 1.71276520685633E-16 ub = 8.232617299999999E-19
+ uc = -8.496648345732E-11 luc = 5.853789657955614E-17 ud = 0
+ up = 0 lp = 1 eu = 1.67
+ vsat = 2.747193515116E5 lvsat = -0.599512211240353 a0 = 1.202162211768
+ la0 = 2.368761249323215E-6 ags = 0.113179367658 lags = 2.192240953832684E-6
+ b0 = 0 b1 = 0 keta = 0.0292908429136
+ lketa = -3.406780567427679E-7 a1 = 0 a2 = 1.201176
+ la2 = -1.61413965952E-6 rdsw = 531.92 rdswmin = 0
+ rdw = 0 rdwmin = 0 rsw = 0
+ rswmin = 0 prwb = -0.32348 prwg = 0.02
+ wr = 1 voff = -0.1979203813256 lvoff = 1.603341065197807E-8
+ voffl = 0 minv = 0 nfactor = 2.52682923776
+ lnfactor = -2.740163486001133E-7 eta0 = 0.08 etab = -0.07
+ dsub = 0.56 cit = 1E-5 cdsc = 0
+ cdscb = 0 cdscd = 0 pclm = -0.48511023428744
+ lpclm = 4.497984479860201E-6 pdiblc1 = 0.39 pdiblc2 = 6.7956520966272E-3
+ lpdiblc2 = -2.541893417244228E-8 pdiblcb = 5.8355983957548E-4 lpdiblcb = -5.450408255827935E-9
+ drout = 0.56 pscbe1 = 6.926355337644E8 lpscbe1 = 431.9830771882613
+ pscbe2 = 1.0062653780232E-8 lpscbe2 = -4.474406435167058E-15 pvag = 0
+ delta = 0.01 fprout = 0 pdits = 0
+ pditsl = 0 pditsd = 0 lambda = 0
+ vtl = 0 lc = 5E-9 xn = 3
+ alpha0 = 1E-10 alpha1 = 1E-10 beta0 = 4.265271567144001
+ lbeta0 = 4.229338067220769E-6 aigbacc = 0.43 bigbacc = 0.054
+ cigbacc = 0.075 nigbacc = 1 aigbinv = 0.35
+ bigbinv = 0.03 cigbinv = 6E-3 eigbinv = 1.1
+ nigbinv = 3 aigc = 0.43 bigc = 0.054
+ cigc = 0.075 aigsd = 0.43 bigsd = 0.054
+ cigsd = 0.075 dlcig = 0 nigc = 1
+ poxedge = 1 pigcd = 1 ntox = 1
+ toxref = 4.23E-9 agidl = 5.43948492672E-11 lagidl = 3.659138390076355E-16
+ bgidl = 1.309797334248E9 lbgidl = -1.246475770293513E3 cgidl = 300
+ egidl = 0.1 noia = 1.2E41 noib = 2E25
+ noic = 0 em = 4.1E7 af = 1
+ ef = 0.88 kf = 0 lintnoi = -6E-8
+ tnoia = 1.5 tnoib = 3.5 ntnoi = 1
+ rnoia = 0.577 rnoib = 0.37 xpart = 0
+ cgso = {5.932020000000001E-11/sw_func_tox_lv_ratio} cgdo = {5.932020000000001E-11/sw_func_tox_lv_ratio} cgbo = {0/sw_func_tox_lv_ratio}
+ ckappas = 0.6 cf = 1.2E-11 clc = 1E-7
+ cle = 0.6 dlc = -2.56E-9 dwc = 0
+ vfbcv = -0.1446893 noff = 4 voffcv = -0.1375
+ acde = 0.552 moin = 14.504 cgsl = {7.513892E-12/sw_func_tox_lv_ratio}
+ cgdl = {7.513892E-12/sw_func_tox_lv_ratio} ijthsrev = 0.1 ijthsfwd = 0.1
+ xjbvs = 1 bvs = 12.8 jss = 2.17E-5
+ jsws = 8.200000000000001E-10 cjs = {7.433E-04*sw_func_psd_nw_cj} mjs = 0.34629
+ mjsws = 0.26859 cjsws = {9.2435E-11*sw_func_psd_nw_cj} cjswgs = {2.4701E-10*sw_func_psd_nw_cj}
+ mjswgs = 0.70393 pbs = 0.6587 pbsws = 0.7418
+ pbswgs = 1.3925 xrcrg1 = 12 xrcrg2 = 1
+ rbpb = 50 rbpd = 50 rbps = 50
+ rbdb = 50 rbsb = 50 gbmin = 1E-12
+ tnom = 30 ute = -0.3030841708 lute = 1.945038289721574E-8
+ kt1 = -0.4308566724 lkt1 = -8.692142066515156E-8 kt1l = 0
+ kt2 = -0.0355619762 lkt2 = -1.924861543977598E-8 ua1 = 2.003584016000001E-9
+ lua1 = 1.669020407943678E-15 ub1 = -6.183355276000001E-19 lub1 = -1.406157764390848E-24
+ uc1 = 1.026796284E-10 luc1 = 1.37766819940032E-16 at = -2.640535588E5
+ lat = 2.118639010102976 prt = 0 njs = 1.2556
+ xtis = 2 tpb = 1.9551E-3 tpbsw = 1.4242E-4
+ tpbswg = 0 tcj = 1.2407E-3 tcjsw = 0
+ tcjswg = 2E-12 tvoff = 0 tvfbsdoff = 0
+ saref = 3E-6 sbref = 3E-6 wlod = 0
+ ku0 = 4.5E-8 kvsat = 0.4 kvth0 = 2.65E-8
+ tku0 = 0 llodku0 = 0 wlodku0 = 1
+ llodvth = 0 wlodvth = 1 lku0 = 0
+ wku0 = 2.5E-7 pku0 = 0 lkvth0 = 0
+ wkvth0 = 2.5E-7 pkvth0 = 0 stk2 = 0
+ lodk2 = 1 steta0 = 0 lodeta0 = 1

.model phighvt_model.3 pmos
+ level = 54 lmin = 2E-6 lmax = 4E-6 wmin = 7E-6
+ wmax = 1.01E-3 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 4.23E-9
+ toxm = 4.23E-9 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 9.999999999999999E22 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {9.364E-9+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {-1.176E-8-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = -5.722E-9 dwb = -1.7864E-8 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = -1.113561301104 lvth0 = 2.85585470499661E-8
+ k1 = 0.3637621455776 lk1 = 2.652566895440147E-7 k2 = 0.05980424599648
+ lk2 = -1.021606893423172E-7 k3 = -13.778 k3b = 2
+ w0 = 0 lpe0 = 0 lpeb = 0
+ vbm = -3 dvtp0 = 0 dvtp1 = 0
+ dvt0 = 4.05 dvt1 = 0.3 dvt2 = 0.03
+ dvt0w = -4.254 dvt1w = 1.1472E6 dvt2w = -8.96E-3
+ vfbsdoff = 0 u0 = 0.014572133174712 lu0 = -9.04081393127723E-9
+ ua = 2.544713549416E-10 lua = -1.896398861498626E-15 ub = 5.914619448359999E-19
+ lub = 9.358961209534573E-25 uc = -6.801805383112002E-11 luc = -9.654448990052035E-18
+ ud = 0 up = 0 lp = 1
+ eu = 1.67 vsat = 1.9525755239136E5 lvsat = -0.279796073244085
+ a0 = 1.862834827728 la0 = -2.894682344441618E-7 ags = 0.4895224060224
+ lags = 6.780172121127532E-7 b0 = 0 b1 = 0
+ keta = -0.05304568723752 lketa = -9.39538094913352E-9 a1 = 0
+ a2 = 0.8 rdsw = 531.92 rdswmin = 0
+ rdw = 0 rdwmin = 0 rsw = 0
+ rswmin = 0 prwb = -0.32348 prwg = 0.02
+ wr = 1 voff = -0.1910957329728 lvoff = -1.142569848847968E-8
+ voffl = 0 minv = 0 nfactor = 2.933877032336
+ lnfactor = -1.911781291032544E-6 eta0 = 0.16043492 leta0 = -3.236315093184E-7
+ etab = -0.14031732 letab = 2.829231433664E-7 dsub = 0.771920062556
+ ldsub = -8.526646100953172E-7 cit = 1E-5 cdsc = 0
+ cdscb = 0 cdscd = 0 pclm = 0.6568215445648
+ lpclm = -9.660087098736425E-8 pdiblc1 = 0.39 pdiblc2 = 7.150215988168E-4
+ lpdiblc2 = -9.533957518921712E-10 pdiblcb = 6.670580670399963E-6 lpdiblcb = -3.129282784838168E-9
+ drout = 0.56 pscbe1 = 8E8 pscbe2 = 9.231951843104E-9
+ lpscbe2 = -1.132060577093806E-15 pvag = 0 delta = 0.01
+ fprout = 0 pdits = 0 pditsl = 0
+ pditsd = 0 lambda = 0 vtl = 0
+ lc = 5E-9 xn = 3 alpha0 = 1E-10
+ alpha1 = 1E-10 beta0 = 3.317690081192 lbeta0 = 8.041951127578366E-6
+ aigbacc = 0.43 bigbacc = 0.054 cigbacc = 0.075
+ nigbacc = 1 aigbinv = 0.35 bigbinv = 0.03
+ cigbinv = 6E-3 eigbinv = 1.1 nigbinv = 3
+ aigc = 0.43 bigc = 0.054 cigc = 0.075
+ aigsd = 0.43 bigsd = 0.054 cigsd = 0.075
+ dlcig = 0 nigc = 1 poxedge = 1
+ pigcd = 1 ntox = 1 toxref = 4.23E-9
+ agidl = 1.858702119504E-10 lagidl = -1.630799122554734E-16 bgidl = 1E9
+ cgidl = 300 egidl = 0.1 noia = 1.2E41
+ noib = 2E25 noic = 0 em = 4.1E7
+ af = 1 ef = 0.88 kf = 0
+ lintnoi = -6E-8 tnoia = 1.5 tnoib = 3.5
+ ntnoi = 1 rnoia = 0.577 rnoib = 0.37
+ xpart = 0 cgso = {5.932020000000001E-11/sw_func_tox_lv_ratio} cgdo = {5.932020000000001E-11/sw_func_tox_lv_ratio}
+ cgbo = {0/sw_func_tox_lv_ratio} ckappas = 0.6 cf = 1.2E-11
+ clc = 1E-7 cle = 0.6 dlc = -2.56E-9
+ dwc = 0 vfbcv = -0.1446893 noff = 4
+ voffcv = -0.1375 acde = 0.552 moin = 14.504
+ cgsl = {7.513892E-12/sw_func_tox_lv_ratio} cgdl = {7.513892E-12/sw_func_tox_lv_ratio} ijthsrev = 0.1
+ ijthsfwd = 0.1 xjbvs = 1 bvs = 12.8
+ jss = 2.17E-5 jsws = 8.200000000000001E-10 cjs = {7.433E-04*sw_func_psd_nw_cj}
+ mjs = 0.34629 mjsws = 0.26859 cjsws = {9.2435E-11*sw_func_psd_nw_cj}
+ cjswgs = {2.4701E-10*sw_func_psd_nw_cj} mjswgs = 0.70393 pbs = 0.6587
+ pbsws = 0.7418 pbswgs = 1.3925 xrcrg1 = 12
+ xrcrg2 = 1 rbpb = 50 rbpd = 50
+ rbps = 50 rbdb = 50 rbsb = 50
+ gbmin = 1E-12 tnom = 30 ute = -0.43143505112
+ lute = 5.358727168823424E-7 kt1 = -0.4745062504 lkt1 = 8.870352940940789E-8
+ kt1l = 0 kt2 = -0.03695862752 lkt2 = -1.362916092072959E-8
+ ua1 = 3.008458432E-9 lua1 = -2.374111902320639E-15 ub1 = -1.3030363232E-18
+ lub1 = 1.348749580721664E-24 uc1 = 3.486156036E-10 luc1 = -8.51761494996672E-16
+ at = 4.361381335999999E5 lat = -0.698596268102272 prt = 0
+ njs = 1.2556 xtis = 2 tpb = 1.9551E-3
+ tpbsw = 1.4242E-4 tpbswg = 0 tcj = 1.2407E-3
+ tcjsw = 0 tcjswg = 2E-12 tvoff = 0
+ tvfbsdoff = 0 saref = 3E-6 sbref = 3E-6
+ wlod = 0 ku0 = 4.5E-8 kvsat = 0.4
+ kvth0 = 2.65E-8 tku0 = 0 llodku0 = 0
+ wlodku0 = 1 llodvth = 0 wlodvth = 1
+ lku0 = 0 wku0 = 2.5E-7 pku0 = 0
+ lkvth0 = 0 wkvth0 = 2.5E-7 pkvth0 = 0
+ stk2 = 0 lodk2 = 1 steta0 = 0
+ lodeta0 = 1

.model phighvt_model.4 pmos
+ level = 54 lmin = 1E-6 lmax = 2E-6 wmin = 7E-6
+ wmax = 1.01E-3 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 4.23E-9
+ toxm = 4.23E-9 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 9.999999999999999E22 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {9.364E-9+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {-1.176E-8-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = -5.722E-9 dwb = -1.7864E-8 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = -1.114072360816 lvth0 = 2.959268659839238E-8
+ k1 = 0.5462826425712 lk1 = -1.040771865324745E-7 k2 = -8.311776183199997E-3
+ lk2 = 3.567344385870886E-8 k3 = -13.778 k3b = 2
+ w0 = 0 lpe0 = 0 lpeb = 0
+ vbm = -3 dvtp0 = 0 dvtp1 = 0
+ dvt0 = 4.05 dvt1 = 0.3 dvt2 = 0.03
+ dvt0w = -4.254 dvt1w = 1.1472E6 dvt2w = -8.96E-3
+ vfbsdoff = 0 u0 = 0.010169809300848 lu0 = -1.326235260359468E-10
+ ua = -7.135920468192E-10 lua = 6.249679323238765E-17 ub = 1.1166695551024E-18
+ lub = -1.268719825728085E-25 uc = -8.182089778416001E-11 luc = 1.827588180580345E-17
+ ud = 0 up = 0 lp = 1
+ eu = 1.67 vsat = 2.447379951472E4 lvsat = 0.065788266376854
+ a0 = 1.7396290528 la0 = -4.015888476185603E-8 ags = 0.6669594002016
+ lags = 3.189699056512583E-7 b0 = 0 b1 = 0
+ keta = -0.07382040309712 lketa = 3.264267208708426E-8 a1 = 0
+ a2 = 0.8 rdsw = 531.92 rdswmin = 0
+ rdw = 0 rdwmin = 0 rsw = 0
+ rswmin = 0 prwb = -0.32348 prwg = 0.02
+ wr = 1 voff = -0.1885326489024 lvoff = -1.661215036661556E-8
+ voffl = 0 minv = 0 nfactor = 2.4768693451664
+ lnfactor = -9.870170958911135E-7 eta0 = -0.2239388882928 leta0 = 4.541565792382466E-7
+ etab = 1.175999999999987E-5 letab = -1.0355565952E-9 dsub = -0.314188925112
+ ldsub = 1.345098648630634E-6 cit = 1E-5 cdsc = 0
+ cdscb = 0 cdscd = 0 pclm = 0.4935007665952
+ lpclm = 2.338819896496808E-7 pdiblc1 = 0.4365156882656 lpdiblc1 = -9.412542551920693E-8
+ pdiblc2 = 5.335115374560003E-5 lpdiblc2 = 3.855076271183034E-10 pdiblcb = -1.744019420784E-3
+ lpdiblcb = 4.132734469048395E-10 drout = 0.2637846837264 ldrout = 5.993976167859548E-7
+ pscbe1 = 8E8 pscbe2 = 8.230625622080002E-9 lpscbe2 = 8.94143057672676E-16
+ pvag = 0 delta = 0.01 fprout = 0
+ pdits = 0 pditsl = 0 pditsd = 0
+ lambda = 0 vtl = 0 lc = 5E-9
+ xn = 3 alpha0 = 1E-10 alpha1 = 1E-10
+ beta0 = 5.736193757504001 lbeta0 = 3.148060568487504E-6 aigbacc = 0.43
+ bigbacc = 0.054 cigbacc = 0.075 nigbacc = 1
+ aigbinv = 0.35 bigbinv = 0.03 cigbinv = 6E-3
+ eigbinv = 1.1 nigbinv = 3 aigc = 0.43
+ bigc = 0.054 cigc = 0.075 aigsd = 0.43
+ bigsd = 0.054 cigsd = 0.075 dlcig = 0
+ nigc = 1 poxedge = 1 pigcd = 1
+ ntox = 1 toxref = 4.23E-9 agidl = 1.106801790304E-10
+ lagidl = -1.093137684119501E-17 bgidl = 8.70486747408E8 lbgidl = 262.0726568849638
+ cgidl = 300 egidl = 0.1 noia = 1.2E41
+ noib = 2E25 noic = 0 em = 4.1E7
+ af = 1 ef = 0.88 kf = 0
+ lintnoi = -6E-8 tnoia = 1.5 tnoib = 3.5
+ ntnoi = 1 rnoia = 0.577 rnoib = 0.37
+ xpart = 0 cgso = {5.932020000000001E-11/sw_func_tox_lv_ratio} cgdo = {5.932020000000001E-11/sw_func_tox_lv_ratio}
+ cgbo = {0/sw_func_tox_lv_ratio} ckappas = 0.6 cf = 1.2E-11
+ clc = 1E-7 cle = 0.6 dlc = -2.56E-9
+ dwc = 0 vfbcv = -0.1446893 noff = 4
+ voffcv = -0.1375 acde = 0.552 moin = 14.504
+ cgsl = {7.513892E-12/sw_func_tox_lv_ratio} cgdl = {7.513892E-12/sw_func_tox_lv_ratio} ijthsrev = 0.1
+ ijthsfwd = 0.1 xjbvs = 1 bvs = 12.8
+ jss = 2.17E-5 jsws = 8.200000000000001E-10 cjs = {7.433E-04*sw_func_psd_nw_cj}
+ mjs = 0.34629 mjsws = 0.26859 cjsws = {9.2435E-11*sw_func_psd_nw_cj}
+ cjswgs = {2.4701E-10*sw_func_psd_nw_cj} mjswgs = 0.70393 pbs = 0.6587
+ pbsws = 0.7418 pbswgs = 1.3925 xrcrg1 = 12
+ xrcrg2 = 1 rbpb = 50 rbpd = 50
+ rbps = 50 rbdb = 50 rbsb = 50
+ gbmin = 1E-12 tnom = 30 ute = 1.106661846912
+ lute = -2.57649711822337E-6 kt1 = -0.3895163794864 lkt1 = -8.327517418167986E-8
+ kt1l = 0 kt2 = -0.04011970337328 lkt2 = -7.232660710100454E-9
+ ua1 = 4.3736668130912E-9 lua1 = -5.136638365626304E-15 ub1 = -2.0702692003824E-18
+ lub1 = 2.901260652357794E-24 uc1 = -1.460855110764704E-10 luc1 = 1.492761045734594E-16
+ at = 3.408125235840002E4 lat = 0.11497387222773 prt = 0
+ njs = 1.2556 xtis = 2 tpb = 1.9551E-3
+ tpbsw = 1.4242E-4 tpbswg = 0 tcj = 1.2407E-3
+ tcjsw = 0 tcjswg = 2E-12 tvoff = 0
+ tvfbsdoff = 0 saref = 3E-6 sbref = 3E-6
+ wlod = 0 ku0 = 4.5E-8 kvsat = 0.4
+ kvth0 = 2.65E-8 tku0 = 0 llodku0 = 0
+ wlodku0 = 1 llodvth = 0 wlodvth = 1
+ lku0 = 0 wku0 = 2.5E-7 pku0 = 0
+ lkvth0 = 0 wkvth0 = 2.5E-7 pkvth0 = 0
+ stk2 = 0 lodk2 = 1 steta0 = 0
+ lodeta0 = 1

.model phighvt_model.5 pmos
+ level = 54 lmin = 5E-7 lmax = 1E-6 wmin = 7E-6
+ wmax = 1.01E-3 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 4.23E-9
+ toxm = 4.23E-9 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 9.999999999999999E22 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {9.364E-9+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {-1.176E-8-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = -5.722E-9 dwb = -1.7864E-8 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = -1.103848212256 lvth0 = 1.912806606426106E-8
+ k1 = 0.4081553230272 lk1 = 3.729888756720023E-8 k2 = 0.03856635403808
+ lk2 = -1.230725998537564E-8 k3 = -13.778 k3b = 2
+ w0 = 0 lpe0 = 0 lpeb = 0
+ vbm = -3 dvtp0 = 0 dvtp1 = 0
+ dvt0 = 4.05 dvt1 = 0.3 dvt2 = 0.03
+ dvt0w = -4.254 dvt1w = 1.1472E6 dvt2w = -8.96E-3
+ vfbsdoff = 0 u0 = 0.012394537811136 lu0 = -2.409677650885917E-9
+ ua = -1.1409003296E-10 lua = -5.511055079927807E-16 ub = 6.999324073311999E-19
+ lub = 2.996668229139702E-25 uc = -1.1534989269216E-10 luc = 5.25934786740396E-17
+ ud = 0 up = 0 lp = 1
+ eu = 1.67 vsat = 6.920653067231999E4 lvsat = 0.020003421382427
+ a0 = 2.34588583072 la0 = -6.606748220985343E-7 ags = 1.0240929258912
+ lags = -4.656340056256098E-8 b0 = 0 b1 = 0
+ keta = -0.05361997634176 lketa = 1.196713129443819E-8 a1 = 0
+ a2 = 0.590592 la2 = 2.1433327616E-7 rdsw = 531.92
+ rdswmin = 0 rdw = 0 rdwmin = 0
+ rsw = 0 rswmin = 0 prwb = -0.32348
+ prwg = 0.02 wr = 1 voff = -0.2184624161856
+ lvoff = 1.40215650430853E-8 voffl = 0 minv = 0
+ nfactor = 0.1665305596512 lnfactor = 1.377660857859404E-6 eta0 = 0.43504927291072
+ leta0 = -2.203309835167801E-7 etab = -1E-3 dsub = 1
+ cit = 1E-5 cdsc = 0 cdscb = 0
+ cdscd = 0 pclm = 0.54700887376 lpclm = 1.791153718043648E-7
+ pdiblc1 = 0.64689936766592 lpdiblc1 = -3.094573290590224E-7 pdiblc2 = 6.70468402944E-5
+ lpdiblc2 = 3.714898180218757E-10 pdiblcb = 0.023432469378688 lpdiblcb = -2.535536636913074E-8
+ drout = 0.7406998475232 ldrout = 1.112654083366544E-7 pscbe1 = 8.42964710528E8
+ lpscbe1 = -43.97524051961856 pscbe2 = 9.071555936672E-9 lpscbe2 = 3.343406208147534E-17
+ pvag = 0 delta = 0.01 fprout = 0
+ pdits = 0 pditsl = 0 pditsd = 0
+ lambda = 0 vtl = 0 lc = 5E-9
+ xn = 3 alpha0 = 1E-10 alpha1 = 1E-10
+ beta0 = 8.54173362784 lbeta0 = 2.765344004012042E-7 aigbacc = 0.43
+ bigbacc = 0.054 cigbacc = 0.075 nigbacc = 1
+ aigbinv = 0.35 bigbinv = 0.03 cigbinv = 6E-3
+ eigbinv = 1.1 nigbinv = 3 aigc = 0.43
+ bigc = 0.054 cigc = 0.075 aigsd = 0.43
+ bigsd = 0.054 cigsd = 0.075 dlcig = 0
+ nigc = 1 poxedge = 1 pigcd = 1
+ ntox = 1 toxref = 4.23E-9 agidl = 1E-10
+ bgidl = 1.081959267296E9 lbgidl = 45.62630332919808 cgidl = 300
+ egidl = 0.1 noia = 1.2E41 noib = 2E25
+ noic = 0 em = 4.1E7 af = 1
+ ef = 0.88 kf = 0 lintnoi = -6E-8
+ tnoia = 1.5 tnoib = 3.5 ntnoi = 1
+ rnoia = 0.577 rnoib = 0.37 xpart = 0
+ cgso = {5.932020000000001E-11/sw_func_tox_lv_ratio} cgdo = {5.932020000000001E-11/sw_func_tox_lv_ratio} cgbo = {0/sw_func_tox_lv_ratio}
+ ckappas = 0.6 cf = 1.2E-11 clc = 1E-7
+ cle = 0.6 dlc = -2.56E-9 dwc = 0
+ vfbcv = -0.1446893 noff = 4 voffcv = -0.1375
+ acde = 0.552 moin = 14.504 cgsl = {7.513892E-12/sw_func_tox_lv_ratio}
+ cgdl = {7.513892E-12/sw_func_tox_lv_ratio} ijthsrev = 0.1 ijthsfwd = 0.1
+ xjbvs = 1 bvs = 12.8 jss = 2.17E-5
+ jsws = 8.200000000000001E-10 cjs = {7.433E-04*sw_func_psd_nw_cj} mjs = 0.34629
+ mjsws = 0.26859 cjsws = {9.2435E-11*sw_func_psd_nw_cj} cjswgs = {2.4701E-10*sw_func_psd_nw_cj}
+ mjswgs = 0.70393 pbs = 0.6587 pbsws = 0.7418
+ pbswgs = 1.3925 xrcrg1 = 12 xrcrg2 = 1
+ rbpb = 50 rbpd = 50 rbps = 50
+ rbdb = 50 rbsb = 50 gbmin = 1E-12
+ tnom = 30 ute = -2.772438769344 lute = 1.393839944526971E-6
+ kt1 = -0.4504618331552 lkt1 = -2.08962834425897E-8 kt1l = 0
+ kt2 = -0.06239031679136 lkt2 = 1.556175753557278E-8 ua1 = -4.0074339781824E-9
+ lua1 = 3.44158591625805E-15 ub1 = 3.7468382087648E-18 lub1 = -3.052665123052548E-24
+ uc1 = 2.040266216537408E-10 luc1 = -2.090706655185664E-16 at = 2.578318312832E5
+ lat = -0.114039320313381 prt = 0 njs = 1.2556
+ xtis = 2 tpb = 1.9551E-3 tpbsw = 1.4242E-4
+ tpbswg = 0 tcj = 1.2407E-3 tcjsw = 0
+ tcjswg = 2E-12 tvoff = 0 tvfbsdoff = 0
+ saref = 2.75E-6 sbref = 2.74E-6 wlod = 0
+ ku0 = 4.5E-8 kvsat = 0.4 kvth0 = 2.65E-8
+ tku0 = 0 llodku0 = 0 wlodku0 = 1
+ llodvth = 0 wlodvth = 1 lku0 = 0
+ wku0 = 2.5E-7 pku0 = 0 lkvth0 = 0
+ wkvth0 = 2.5E-7 pkvth0 = 0 stk2 = 0
+ lodk2 = 1 steta0 = 0 lodeta0 = 1

.model phighvt_model.6 pmos
+ level = 54 lmin = 2.5E-7 lmax = 5E-7 wmin = 7E-6
+ wmax = 1.01E-3 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 4.23E-9
+ toxm = 4.23E-9 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 9.999999999999999E22 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {9.364E-9+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {-1.176E-8-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = -5.722E-9 dwb = -1.7864E-8 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = -1.074569583168 lvth0 = 3.800118164111322E-9
+ k1 = 0.1864214550336 lk1 = 1.533810021392097E-7 k2 = 0.11639874788736
+ lk2 = -5.30540748133507E-8 k3 = -13.778 k3b = 2
+ w0 = 0 lpe0 = 0 lpeb = 0
+ vbm = -3 dvtp0 = 0 dvtp1 = 0
+ dvt0 = 4.05 dvt1 = 0.3 dvt2 = 0.03
+ dvt0w = -4.254 dvt1w = 1.1472E6 dvt2w = -8.96E-3
+ vfbsdoff = 0 u0 = 0.0110571021088 lu0 = -1.709503311998976E-9
+ ua = -3.892222603839998E-10 lua = -4.070682842917683E-16 ub = 8.021372384000003E-19
+ lub = 2.461605497528319E-25 uc = -3.120030036410848E-11 luc = 8.539484098458069E-18
+ ud = 0 up = 0 lp = 1
+ eu = 1.67 vsat = 1.345026856E5 lvsat = -0.014180421645312
+ a0 = 1.414257456 la0 = -1.7294873536512E-7 ags = -0.564888384
+ lags = 7.853000947916798E-7 b0 = 0 b1 = 0
+ keta = 0.03131491104 lketa = -3.249798094766079E-8 a1 = 0
+ a2 = 1.218816 la2 = -1.1455455232E-7 rdsw = 531.92
+ rdswmin = 0 rdw = 0 rdwmin = 0
+ rsw = 0 rswmin = 0 prwb = -0.32348
+ prwg = 0.02 wr = 1 voff = -0.1541734073888
+ lvoff = -1.963501684221542E-8 voffl = 0 minv = 0
+ nfactor = 3.758949631456 lnfactor = -5.03042374611845E-7 eta0 = -0.50639515265024
+ leta0 = 2.725340021528936E-7 etab = -1.41028E-3 letab = 2.147897856E-10
+ dsub = 1.346256134224 ldsub = -1.812720113889484E-7 cit = 1E-5
+ cdsc = 0 cdscb = 0 cdscd = 0
+ pclm = 1.071829846224 lpclm = -9.563890369998843E-8 pdiblc1 = -0.29324550944064
+ lpdiblc1 = 1.827273170038038E-7 pdiblc2 = -7.641251795788799E-3 lpdiblc2 = 4.406938319984152E-9
+ pdiblcb = -0.025 drout = 1.3811077335136 ldrout = -2.240009281370399E-7
+ pscbe1 = 7.14070578944E8 lpscbe1 = 23.503415247237115 pscbe2 = 1.8036220104192E-8
+ lpscbe2 = -4.659746922898595E-15 pvag = 0 delta = 0.01
+ fprout = 0 pdits = 0 pditsl = 0
+ pditsd = 0 lambda = 0 vtl = 0
+ lc = 5E-9 xn = 3 alpha0 = -1.705613500224E-8
+ lalpha0 = 8.981579796372685E-15 alpha1 = 2.09408E-10 lalpha1 = -5.727727616E-17
+ beta0 = 0.777889648192002 lbeta0 = 4.341062000626523E-6 aigbacc = 0.43
+ bigbacc = 0.054 cigbacc = 0.075 nigbacc = 1
+ aigbinv = 0.35 bigbinv = 0.03 cigbinv = 6E-3
+ eigbinv = 1.1 nigbinv = 3 aigc = 0.43
+ bigc = 0.054 cigc = 0.075 aigsd = 0.43
+ bigsd = 0.054 cigsd = 0.075 dlcig = 0
+ nigc = 1 poxedge = 1 pigcd = 1
+ ntox = 1 toxref = 4.23E-9 agidl = 1E-10
+ bgidl = 1.089046440928E9 lbgidl = 41.91602618937343 cgidl = 300
+ egidl = 0.1 noia = 1.2E41 noib = 2E25
+ noic = 0 em = 4.1E7 af = 1
+ ef = 0.88 kf = 0 lintnoi = -6E-8
+ tnoia = 1.5 tnoib = 3.5 ntnoi = 1
+ rnoia = 0.577 rnoib = 0.37 xpart = 0
+ cgso = {5.932020000000001E-11/sw_func_tox_lv_ratio} cgdo = {5.932020000000001E-11/sw_func_tox_lv_ratio} cgbo = {0/sw_func_tox_lv_ratio}
+ ckappas = 0.6 cf = 1.2E-11 clc = 1E-7
+ cle = 0.6 dlc = -2.56E-9 dwc = 0
+ vfbcv = -0.1446893 noff = 4 voffcv = -0.1375
+ acde = 0.552 moin = 14.504 cgsl = {7.513892E-12/sw_func_tox_lv_ratio}
+ cgdl = {7.513892E-12/sw_func_tox_lv_ratio} ijthsrev = 0.1 ijthsfwd = 0.1
+ xjbvs = 1 bvs = 12.8 jss = 2.17E-5
+ jsws = 8.200000000000001E-10 cjs = {7.433E-04*sw_func_psd_nw_cj} mjs = 0.34629
+ mjsws = 0.26859 cjsws = {9.2435E-11*sw_func_psd_nw_cj} cjswgs = {2.4701E-10*sw_func_psd_nw_cj}
+ mjswgs = 0.70393 pbs = 0.6587 pbsws = 0.7418
+ pbswgs = 1.3925 xrcrg1 = 12 xrcrg2 = 1
+ rbpb = 50 rbpd = 50 rbps = 50
+ rbdb = 50 rbsb = 50 gbmin = 1E-12
+ tnom = 30 ute = -0.1756448 lute = 3.4366365696E-8
+ kt1 = -0.4832542079104 lkt1 = -3.728819410747396E-9 kt1l = 0
+ kt2 = -0.026421654776 lkt2 = -3.268556402708478E-9 ua1 = 4.058230268704E-9
+ lua1 = -7.809506302719181E-16 ub1 = -3.5516770096064E-18 lub1 = 7.682535640691424E-25
+ uc1 = -3.279197338524799E-10 luc1 = 6.941389051605031E-17 at = 3.421565593216001E4
+ lat = 3.028219806395594E-3 prt = 0 njs = 1.2556
+ xtis = 2 tpb = 1.9551E-3 tpbsw = 1.4242E-4
+ tpbswg = 0 tcj = 1.2407E-3 tcjsw = 0
+ tcjswg = 2E-12 tvoff = 0 tvfbsdoff = 0
+ saref = 1.75E-6 sbref = 1.74E-6 wlod = 0
+ ku0 = 4.5E-8 kvsat = 0.4 kvth0 = 2.65E-8
+ tku0 = 0 llodku0 = 0 wlodku0 = 1
+ llodvth = 0 wlodvth = 1 lku0 = 0
+ wku0 = 2.5E-7 pku0 = 0 lkvth0 = 0
+ wkvth0 = 2.5E-7 pkvth0 = 0 stk2 = 0
+ lodk2 = 1 steta0 = 0 lodeta0 = 1

.model phighvt_model.7 pmos
+ level = 54 lmin = 1.8E-7 lmax = 2.5E-7 wmin = 7E-6
+ wmax = 1.01E-3 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 4.23E-9
+ toxm = 4.23E-9 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 9.999999999999999E22 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {9.364E-9+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {-1.176E-8-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = -5.722E-9 dwb = -1.7864E-8 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = -0.993875702628572 lvth0 = -1.827127204103315E-8
+ k1 = 0.058378083725714 lk1 = 1.884034250593427E-7 k2 = 0.192597518102857
+ lk2 = -7.389596244269353E-8 k3 = -13.778 k3b = 2
+ w0 = 0 lpe0 = 0 lpeb = 0
+ vbm = -3 dvtp0 = 0 dvtp1 = 0
+ dvt0 = 4.05 dvt1 = 0.3 dvt2 = 0.03
+ dvt0w = -4.254 dvt1w = 1.1472E6 dvt2w = -8.96E-3
+ vfbsdoff = 0 u0 = 8.955263714285719E-3 lu0 = -1.134608474331429E-9
+ ua = -6.936577566857133E-10 lua = -3.237990873433237E-16 ub = 8.830292228571413E-19
+ lub = 2.240349741641147E-25 uc = 3.188619753810174E-11 luc = -8.715934807754466E-18
+ ud = 0 up = 0 lp = 1
+ eu = 1.67 vsat = 3.441989885714282E4 lvsat = 0.013194222184594
+ a0 = 1.296564857142858 la0 = -1.407574557257144E-7 ags = 5.37702605714286
+ lags = -8.399323431497149E-7 b0 = 0 b1 = 0
+ keta = -0.085414373714286 lketa = -5.701869816685792E-10 a1 = 0
+ a2 = 1.019254421942857 la2 = -5.997046948981035E-8 rdsw = 531.92
+ rdswmin = 0 rdw = 0 rdwmin = 0
+ rsw = 0 rswmin = 0 prwb = -0.32348
+ prwg = 0.02 wr = 1 voff = -0.138161020331429
+ lvoff = -2.401472495014766E-8 voffl = 0 minv = 0
+ nfactor = 2.282860503885715 lnfactor = -9.930247643882064E-8 eta0 = 0.49
+ etab = -6.25E-4 dsub = 1.028118281405715 ldsub = -9.425494588609103E-8
+ cit = 1E-5 cdsc = 0 cdscb = 0
+ cdscd = 0 pclm = 0.777310028971429 lpclm = -1.508184328506514E-8
+ pdiblc1 = 0.279541629085714 lpdiblc1 = 2.605857887407547E-8 pdiblc2 = 6.534625464228569E-3
+ lpdiblc2 = 5.295523718242016E-10 pdiblcb = 0.412248967862858 lpdiblcb = -1.195963376898488E-7
+ drout = 0.495473916857143 ldrout = 1.823763339483425E-8 pscbe1 = 8E8
+ pscbe2 = -2.307990462354287E-8 lpscbe2 = 6.586335512631446E-15 pvag = 0
+ delta = 0.01 fprout = 0 pdits = 0
+ pditsl = 0 pditsd = 0 lambda = 0
+ vtl = 0 lc = 5E-9 xn = 3
+ alpha0 = 1.947043974628572E-8 lalpha0 = -1.009168928844071E-15 alpha1 = 0
+ beta0 = 17.99855519428571 lbeta0 = -3.69134439541028E-7 aigbacc = 0.43
+ bigbacc = 0.054 cigbacc = 0.075 nigbacc = 1
+ aigbinv = 0.35 bigbinv = 0.03 cigbinv = 6E-3
+ eigbinv = 1.1 nigbinv = 3 aigc = 0.43
+ bigc = 0.054 cigc = 0.075 aigsd = 0.43
+ bigsd = 0.054 cigsd = 0.075 dlcig = 0
+ nigc = 1 poxedge = 1 pigcd = 1
+ ntox = 1 toxref = 4.23E-9 agidl = 1E-10
+ bgidl = 7.917466295999997E8 lbgidl = 123.23347058380809 cgidl = 1.029648303360001E3
+ lcgidl = -1.995734039350273E-4 egidl = 0.1 noia = 1.2E41
+ noib = 2E25 noic = 0 em = 4.1E7
+ af = 1 ef = 0.88 kf = 0
+ lintnoi = -6E-8 tnoia = 1.5 tnoib = 3.5
+ ntnoi = 1 rnoia = 0.577 rnoib = 0.37
+ xpart = 0 cgso = {5.932020000000001E-11/sw_func_tox_lv_ratio} cgdo = {5.932020000000001E-11/sw_func_tox_lv_ratio}
+ cgbo = {0/sw_func_tox_lv_ratio} ckappas = 0.6 cf = 1.2E-11
+ clc = 1E-7 cle = 0.6 dlc = -2.56E-9
+ dwc = 0 vfbcv = -0.1446893 noff = 4
+ voffcv = -0.1375 acde = 0.552 moin = 14.504
+ cgsl = {7.513892E-12/sw_func_tox_lv_ratio} cgdl = {7.513892E-12/sw_func_tox_lv_ratio} ijthsrev = 0.1
+ ijthsfwd = 0.1 xjbvs = 1 bvs = 12.8
+ jss = 2.17E-5 jsws = 8.200000000000001E-10 cjs = {7.433E-04*sw_func_psd_nw_cj}
+ mjs = 0.34629 mjsws = 0.26859 cjsws = {9.2435E-11*sw_func_psd_nw_cj}
+ cjswgs = {2.4701E-10*sw_func_psd_nw_cj} mjswgs = 0.70393 pbs = 0.6587
+ pbsws = 0.7418 pbswgs = 1.3925 xrcrg1 = 12
+ xrcrg2 = 1 rbpb = 50 rbpd = 50
+ rbps = 50 rbdb = 50 rbsb = 50
+ gbmin = 1E-12 tnom = 30 ute = 0.289994697142857
+ lute = -9.299534956251434E-8 kt1 = -0.436403450834286 lkt1 = -1.654343848620616E-8
+ kt1l = 0 kt2 = 4.409361470857187E-3 lkt2 = -1.170145596654886E-8
+ ua1 = 3.602933223200002E-9 lua1 = -6.564177823856644E-16 ub1 = -3.107637687977145E-18
+ lub1 = 6.467999288171086E-25 uc1 = -2.624919929040002E-10 luc1 = 5.151809481182211E-17
+ at = 8.092896367085716E4 lat = -9.74880412629285E-3 prt = 0
+ njs = 1.2556 xtis = 2 tpb = 1.9551E-3
+ tpbsw = 1.4242E-4 tpbswg = 0 tcj = 1.2407E-3
+ tcjsw = 0 tcjswg = 2E-12 tvoff = 0
+ tvfbsdoff = 0 saref = 1.25E-6 sbref = 1.24E-6
+ wlod = 0 ku0 = 4.5E-8 kvsat = 0.4
+ kvth0 = 2.65E-8 tku0 = 0 llodku0 = 0
+ wlodku0 = 1 llodvth = 0 wlodvth = 1
+ lku0 = 0 wku0 = 2.5E-7 pku0 = 0
+ lkvth0 = 0 wkvth0 = 2.5E-7 pkvth0 = 0
+ stk2 = 0 lodk2 = 1 steta0 = 0
+ lodeta0 = 1

.model phighvt_model.8 pmos
+ level = 54 lmin = 1.5E-7 lmax = 1.8E-7 wmin = 7E-6
+ wmax = 1.01E-3 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 4.23E-9
+ toxm = 4.23E-9 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 9.999999999999999E22 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {9.364E-9+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {-1.176E-8-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = -5.722E-9 dwb = -1.7864E-8 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = -0.958775439999972 lvth0 = -2.54148774912057E-8
+ k1 = 1.750243002399999 lk1 = -1.559249231892477E-7 k2 = -0.570215021279999
+ lk2 = 8.135164557250545E-8 k3 = -13.778 k3b = 2
+ w0 = 0 lpe0 = 0 lpeb = 0
+ vbm = -3 dvtp0 = 0 dvtp1 = 0
+ dvt0 = 4.05 dvt1 = 0.3 dvt2 = 0.03
+ dvt0w = -4.254 dvt1w = 1.1472E6 dvt2w = -8.96E-3
+ vfbsdoff = 0 u0 = 0.01099341432 lu0 = -1.549412885606397E-9
+ ua = -2.31439860800004E-10 lua = -4.178696735139832E-16 ub = 3.700997840000036E-19
+ lub = 3.284263735603193E-25 uc = -1.277637053039998E-10 luc = 2.377601341867004E-17
+ ud = 0 up = 0 lp = 1
+ eu = 1.67 vsat = 2.265384879999998E5 lvsat = -0.02590575307776
+ a0 = -2.641985159999994 la0 = 6.608162437631989E-7 ags = 1.25
+ b0 = 0 b1 = 0 keta = -0.0476400357712
+ lketa = -8.258020239845358E-9 a1 = 0 a2 = 2.298369773999998
+ la2 = -3.202960259404795E-7 rdsw = 531.92 rdswmin = 0
+ rdw = 0 rdwmin = 0 rsw = 0
+ rswmin = 0 prwb = -0.32348 prwg = 0.02
+ wr = 1 voff = -0.22689045512 lvoff = -5.956510381977622E-9
+ voffl = 0 minv = 0 nfactor = 1.056753756800002
+ lnfactor = 1.502347687280637E-7 eta0 = 0.49 etab = -4.203850203519994E-3
+ letab = 7.283675873147892E-10 dsub = 3.130060560000647E-3 ldsub = 1.143506568204287E-7
+ cit = 1E-5 cdsc = 0 cdscb = 0
+ cdscd = 0 pclm = -0.010854379839998 lpclm = 1.453253771962365E-7
+ pdiblc1 = 1.678979306319998 lpdiblc1 = -2.58754977196646E-7 pdiblc2 = -0.1471078324488
+ lpdiblc2 = 3.179886540628371E-8 pdiblcb = 0.11155240832 lpdiblcb = -5.839857389168632E-8
+ drout = -1.803819106079996 ldrout = 4.861897494230008E-7 pscbe1 = 7.9989774E8
+ pscbe2 = 9.078126498399995E-9 lpscbe2 = 4.153301869363271E-17 pvag = 0
+ delta = 0.01 fprout = 0 pdits = 0
+ pditsl = 0 pditsd = 0 lambda = 0
+ vtl = 0 lc = 5E-9 xn = 3
+ alpha0 = 9.787009894399984E-8 lalpha0 = -1.696506756876285E-14 alpha1 = -5.78399999999999E-10
+ lalpha1 = 1.177159679999998E-16 beta0 = 57.248836451999935 lbeta0 = -8.357351681111028E-6
+ aigbacc = 0.43 bigbacc = 0.054 cigbacc = 0.075
+ nigbacc = 1 aigbinv = 0.35 bigbinv = 0.03
+ cigbinv = 6E-3 eigbinv = 1.1 nigbinv = 3
+ aigc = 0.43 bigc = 0.054 cigc = 0.075
+ aigsd = 0.43 bigsd = 0.054 cigsd = 0.075
+ dlcig = 0 nigc = 1 poxedge = 1
+ pigcd = 1 ntox = 1 toxref = 4.23E-9
+ agidl = 4.10752340799999E-10 lagidl = -6.324431639961581E-17 bgidl = 3.694991487999996E9
+ lbgidl = -467.6349229977592 cgidl = -1.402512707839997E3 lcgidl = 2.954200050643963E-4
+ egidl = 0.1 noia = 1.2E41 noib = 2E25
+ noic = 0 em = 4.1E7 af = 1
+ ef = 0.88 kf = 0 lintnoi = -6E-8
+ tnoia = 1.5 tnoib = 3.5 ntnoi = 1
+ rnoia = 0.577 rnoib = 0.37 xpart = 0
+ cgso = {5.932020000000001E-11/sw_func_tox_lv_ratio} cgdo = {5.932020000000001E-11/sw_func_tox_lv_ratio} cgbo = {0/sw_func_tox_lv_ratio}
+ ckappas = 0.6 cf = 1.2E-11 clc = 1E-7
+ cle = 0.6 dlc = -2.56E-9 dwc = 0
+ vfbcv = -0.1446893 noff = 4 voffcv = -0.1375
+ acde = 0.552 moin = 14.504 cgsl = {7.513892E-12/sw_func_tox_lv_ratio}
+ cgdl = {7.513892E-12/sw_func_tox_lv_ratio} ijthsrev = 0.1 ijthsfwd = 0.1
+ xjbvs = 1 bvs = 12.8 jss = 2.17E-5
+ jsws = 8.200000000000001E-10 cjs = {7.433E-04*sw_func_psd_nw_cj} mjs = 0.34629
+ mjsws = 0.26859 cjsws = {9.2435E-11*sw_func_psd_nw_cj} cjswgs = {2.4701E-10*sw_func_psd_nw_cj}
+ mjswgs = 0.70393 pbs = 0.6587 pbsws = 0.7418
+ pbswgs = 1.3925 xrcrg1 = 12 xrcrg2 = 1
+ rbpb = 50 rbpd = 50 rbps = 50
+ rbdb = 50 rbsb = 50 gbmin = 1E-12
+ tnom = 30 ute = -1.002294199999999 lute = 1.700112867839997E-7
+ kt1 = -0.035130880000001 lkt1 = -9.821043210239983E-8 kt1l = 0
+ kt2 = -0.115281352 lkt2 = 1.265799803903998E-8 ua1 = 8.65085519999999E-10
+ lua1 = -9.921101783039981E-17 ub1 = 1.621275359999998E-19 lub1 = -1.866268956671996E-26
+ uc1 = 2.739337871999995E-10 luc1 = -5.76552799549439E-17 at = -9.429519199999976E4
+ lat = 0.02591281603584 prt = 0 njs = 1.2556
+ xtis = 2 tpb = 1.9551E-3 tpbsw = 1.4242E-4
+ tpbswg = 0 tcj = 1.2407E-3 tcjsw = 0
+ tcjswg = 2E-12 tvoff = 0 tvfbsdoff = 0
+ saref = 1.1E-6 sbref = 1.1E-6 wlod = 0
+ ku0 = 4.5E-8 kvsat = 0.4 kvth0 = 2.65E-8
+ tku0 = 0 llodku0 = 0 wlodku0 = 1
+ llodvth = 0 wlodvth = 1 lku0 = 0
+ wku0 = 2.5E-7 pku0 = 0 lkvth0 = 0
+ wkvth0 = 2.5E-7 pkvth0 = 0 stk2 = 0
+ lodk2 = 1 steta0 = 0 lodeta0 = 1

.model phighvt_model.9 pmos
+ level = 54 lmin = 8E-6 lmax = 2.02E-5 wmin = 5E-6
+ wmax = 7E-6 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 4.23E-9
+ toxm = 4.23E-9 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 9.999999999999999E22 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {9.364E-9+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {-1.176E-8-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = -5.722E-9 dwb = -1.7864E-8 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = -1.14246178619 wvth0 = 1.93048131314234E-7
+ k1 = 0.44253196176072 wk1 = -4.160937079014565E-8 k2 = 0.01988271752902
+ wk2 = 7.022161638907954E-8 k3 = -13.778 k3b = 2
+ w0 = 0 lpe0 = 0 lpeb = 0
+ vbm = -3 dvtp0 = 0 dvtp1 = 0
+ dvt0 = 4.05 dvt1 = 0.3 dvt2 = 0.03
+ dvt0w = -4.254 dvt1w = 1.1472E6 dvt2w = -8.96E-3
+ vfbsdoff = 0 u0 = 0.019609501613512 wu0 = -5.227369558131013E-8
+ ua = 1.22586952380964E-9 wua = -1.022022262927542E-14 ub = 1.817906574156796E-19
+ wub = 4.478284037842883E-24 uc = -7.297295053033202E-11 wuc = -3.279623891051997E-17
+ ud = 0 up = 0 lp = 1
+ eu = 1.67 vsat = 2.9884711625E5 wvsat = -0.69007860495687
+ a0 = 1.0040103484704 wa0 = 3.444413357830154E-6 ags = 3.808545616159842E-3
+ wags = 2.671018291815581E-6 b0 = 0 b1 = 0
+ keta = 0.078791664811056 wketa = -6.420029868111146E-7 a1 = 0
+ a2 = 1.4981272 wa2 = -3.4775614737984E-6 rdsw = 531.92
+ rdswmin = 0 rdw = 0 rdwmin = 0
+ rsw = 0 rswmin = 0 prwb = -0.32348
+ prwg = 0.02 wr = 1 voff = -0.09816566306712
+ wvoff = -6.824641363538412E-7 voffl = 0 minv = 0
+ nfactor = 6.5731323865024 wnfactor = -2.848676474827518E-5 eta0 = 0.08
+ etab = -0.07 dsub = 0.56 cit = 1E-5
+ cdsc = 0 cdscb = 0 cdscd = 0
+ pclm = -0.173499662253208 wpclm = 1.738262197707842E-6 pdiblc1 = 0.39
+ pdiblc2 = 0.012248218710457 wpdiblc2 = -6.018288821475584E-8 pdiblcb = 7.300287385315997E-3
+ wpdiblcb = -5.163370709369739E-8 drout = 0.56 pscbe1 = 8.1554559699016E8
+ wpscbe1 = -482.1997172253283 pscbe2 = 9.256113705191204E-9 wpscbe2 = 1.737490561592399E-15
+ pvag = 0 delta = 0.01 fprout = 0
+ pdits = 0 pditsl = 0 pditsd = 0
+ lambda = 0 vtl = 0 lc = 5E-9
+ xn = 3 alpha0 = -8.328613626781999E-10 walpha0 = 6.512558911147163E-15
+ alpha1 = 3.483780042970061E-10 walpha1 = -1.733994406814569E-15 beta0 = 8.7216333899248
+ wbeta0 = -2.74311231424119E-5 aigbacc = 0.43 bigbacc = 0.054
+ cigbacc = 0.075 nigbacc = 1 aigbinv = 0.35
+ bigbinv = 0.03 cigbinv = 6E-3 eigbinv = 1.1
+ nigbinv = 3 aigc = 0.43 bigc = 0.054
+ cigc = 0.075 aigsd = 0.43 bigsd = 0.054
+ cigsd = 0.075 dlcig = 0 nigc = 1
+ poxedge = 1 pigcd = 1 ntox = 1
+ toxref = 4.23E-9 agidl = 1E-10 bgidl = 4.173042634508001E8
+ wbgidl = 5.146177191621507E3 cgidl = 300 egidl = 0.1
+ noia = 1.2E41 noib = 2E25 noic = 0
+ em = 4.1E7 af = 1 ef = 0.88
+ kf = 0 lintnoi = -6E-8 tnoia = 1.5
+ tnoib = 3.5 ntnoi = 1 rnoia = 0.577
+ rnoib = 0.37 xpart = 0 cgso = {5.932020000000001E-11/sw_func_tox_lv_ratio}
+ cgdo = {5.932020000000001E-11/sw_func_tox_lv_ratio} cgbo = {0/sw_func_tox_lv_ratio} ckappas = 0.6
+ cf = 1.2E-11 clc = 1E-7 cle = 0.6
+ dlc = -2.56E-9 dwc = 0 vfbcv = -0.1446893
+ noff = 4 voffcv = -0.1375 acde = 0.552
+ moin = 14.504 cgsl = {7.513892E-12/sw_func_tox_lv_ratio} cgdl = {7.513892E-12/sw_func_tox_lv_ratio}
+ ijthsrev = 0.1 ijthsfwd = 0.1 xjbvs = 1
+ bvs = 12.8 jss = 2.17E-5 jsws = 8.200000000000001E-10
+ cjs = {7.433E-04*sw_func_psd_nw_cj} mjs = 0.34629 mjsws = 0.26859
+ cjsws = {9.2435E-11*sw_func_psd_nw_cj} cjswgs = {2.4701E-10*sw_func_psd_nw_cj} mjswgs = 0.70393
+ pbs = 0.6587 pbsws = 0.7418 pbswgs = 1.3925
+ xrcrg1 = 12 xrcrg2 = 1 rbpb = 50
+ rbpd = 50 rbps = 50 rbdb = 50
+ rbsb = 50 gbmin = 1E-12 tnom = 30
+ ute = -0.17595385548 wute = -8.706075149654295E-7 kt1 = -0.46659636
+ wkt1 = 1.738780736899202E-7 kt1l = 0 kt2 = -0.037961
+ ua1 = 2.2116E-9 ub1 = -4.7735394708E-19 wub1 = -2.207729901640914E-24
+ uc1 = 1.1985E-10 at = 0 prt = 0
+ njs = 1.2556 xtis = 2 tpb = 1.9551E-3
+ tpbsw = 1.4242E-4 tpbswg = 0 tcj = 1.2407E-3
+ tcjsw = 0 tcjswg = 2E-12 tvoff = 0
+ tvfbsdoff = 0 saref = 3E-6 sbref = 3E-6
+ wlod = 0 ku0 = 4.5E-8 kvsat = 0.4
+ kvth0 = 2.65E-8 tku0 = 0 llodku0 = 0
+ wlodku0 = 1 llodvth = 0 wlodvth = 1
+ lku0 = 0 wku0 = 2.5E-7 pku0 = 0
+ lkvth0 = 0 wkvth0 = 2.5E-7 pkvth0 = 0
+ stk2 = 0 lodk2 = 1 steta0 = 0
+ lodeta0 = 1

.model phighvt_model.10 pmos
+ level = 54 lmin = 4E-6 lmax = 8E-6 wmin = 5E-6
+ wmax = 7E-6 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 4.23E-9
+ toxm = 4.23E-9 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 9.999999999999999E22 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {9.364E-9+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {-1.176E-8-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = -5.722E-9 dwb = -1.7864E-8 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = -1.16187819316784 lvth0 = 1.557879297148397E-7
+ wvth0 = 2.699903490519071E-7 pvth0 = -6.173474228625756E-13 k1 = 0.614477387961447
+ lk1 = -1.379607566030056E-6 wk1 = -1.19367146540943E-6 pk1 = 9.24359325741972E-12
+ k2 = -0.056217310596584 lk2 = 6.105900976663468E-7 wk2 = 5.70092198622036E-7
+ pk2 = -4.010721613957771E-12 k3 = -13.778 k3b = 2
+ w0 = 0 lpe0 = 0 lpeb = 0
+ vbm = -3 dvtp0 = 0 dvtp1 = 0
+ dvt0 = 4.05 dvt1 = 0.3 dvt2 = 0.03
+ dvt0w = -4.254 dvt1w = 1.1472E6 dvt2w = -8.96E-3
+ vfbsdoff = 0 u0 = 0.022414066662262 lu0 = -2.250248375994708E-8
+ wu0 = -7.328107404856414E-8 pu0 = 1.68553121279582E-13 ua = 1.894261785275956E-9
+ lua = -5.362858677720214E-15 wua = -1.50354786646371E-14 pua = 3.86353031048452E-20
+ ub = -1.720579304718514E-19 lub = 2.839111221887364E-24 wub = 6.942933633659501E-24
+ pub = -1.977516532502656E-29 uc = -1.288959178455996E-10 luc = 4.486990467133956E-16
+ wuc = 3.066833302707334E-16 puc = -2.72382111291717E-21 ud = 0
+ up = 0 lp = 1 eu = 1.67
+ vsat = 3.971096975806673E5 lvsat = -0.788411786558236 wvsat = -0.85444029608229
+ pvsat = 1.318759315978629E-6 a0 = 0.095306498583764 la0 = 7.291003513642422E-6
+ wa0 = 7.727260798493138E-6 pa0 = -3.436351209710828E-11 ags = -0.660742793711715
+ lags = 5.332040962123994E-6 wags = 5.402961115349877E-6 pags = -2.191979788348389E-11
+ b0 = 0 b1 = 0 keta = 0.223254210910808
+ lketa = -1.159098127882279E-6 wketa = -1.354111030024602E-6 pketa = 5.713613126884278E-12
+ a1 = 0 a2 = 2.200359387936 la2 = -5.634374004548253E-6
+ wa2 = -6.975571009062733E-6 pa2 = 2.806634946638409E-11 rdsw = 531.92
+ rdswmin = 0 rdw = 0 rdwmin = 0
+ rsw = 0 rswmin = 0 prwb = -0.32348
+ prwg = 0.02 wr = 1 voff = -0.059373882033988
+ lvoff = -3.112466309549513E-7 wvoff = -9.672307962025473E-7 pvoff = 2.284830990629292E-12
+ voffl = 0 minv = 0 nfactor = 7.767593116654776
+ lnfactor = -9.583779557592181E-6 wnfactor = -3.658719812633949E-5 pnfactor = 6.499398921756649E-11
+ eta0 = 0.08 etab = -0.07 dsub = 0.56
+ cit = 1E-5 cdsc = 0 cdscb = 0
+ cdscd = 0 pclm = -0.984552940020465 lpclm = 6.50750219523114E-6
+ wpclm = 3.486745377138207E-6 ppclm = -1.402898975982312E-11 pdiblc1 = 0.39
+ pdiblc2 = 0.023428525823621 lpdiblc2 = -8.970541772860968E-8 wpdiblc2 = -1.161186156297971E-7
+ ppdiblc2 = 4.48801427629132E-13 pdiblcb = 9.707473308947818E-3 lpdiblcb = -1.93141044019784E-8
+ wpdiblcb = -6.369652163415197E-8 ppdiblcb = 9.678623372162817E-14 drout = 0.56
+ pscbe1 = 6.407730834590788E8 lpscbe1 = 1.402290757766901E3 wpscbe1 = 362.0658721679304
+ ppscbe1 = -6.7739818418086E-3 pscbe2 = 9.820213557438182E-9 lpscbe2 = -4.526066446500677E-15
+ wpscbe2 = 1.692541139064247E-15 ppscbe2 = 3.606525906430824E-22 pvag = 0
+ delta = 0.01 fprout = 0 pdits = 0
+ pditsl = 0 pditsd = 0 lambda = 0
+ vtl = 0 lc = 5E-9 xn = 3
+ alpha0 = -1.771207950168948E-9 lalpha0 = 7.528842611663765E-15 walpha0 = 1.306341166869187E-14
+ palpha0 = -5.256089811721512E-20 alpha1 = 5.982164712592786E-10 lalpha1 = -2.004583936441132E-15
+ walpha1 = -3.478184700741207E-15 palpha1 = 1.399454570712626E-20 beta0 = 13.780495673216382
+ lbeta0 = -4.058988270723569E-5 wbeta0 = -6.642836762544817E-5 pbeta0 = 3.128951710545312E-10
+ aigbacc = 0.43 bigbacc = 0.054 cigbacc = 0.075
+ nigbacc = 1 aigbinv = 0.35 bigbinv = 0.03
+ cigbinv = 6E-3 eigbinv = 1.1 nigbinv = 3
+ aigc = 0.43 bigc = 0.054 cigc = 0.075
+ aigsd = 0.43 bigsd = 0.054 cigsd = 0.075
+ dlcig = 0 nigc = 1 poxedge = 1
+ pigcd = 1 ntox = 1 toxref = 4.23E-9
+ agidl = 9.321422381096217E-9 lagidl = -7.398826690317314E-14 wagidl = -6.469563983118704E-14
+ pagidl = 5.190867600983259E-19 bgidl = 2.404173694135516E9 lbgidl = -1.594168661448743E4
+ wbgidl = -7.640139038744638E3 pbgidl = 0.102591264000667 cgidl = 300
+ egidl = 0.625564299150895 legidl = -4.216875665523186E-6 wegidl = -3.669107325861765E-6
+ pegidl = 2.943915601119839E-11 noia = 1.2E41 noib = 2E25
+ noic = 0 em = 4.1E7 af = 1
+ ef = 0.88 kf = 0 lintnoi = -6E-8
+ tnoia = 1.5 tnoib = 3.5 ntnoi = 1
+ rnoia = 0.577 rnoib = 0.37 xpart = 0
+ cgso = {5.932020000000001E-11/sw_func_tox_lv_ratio} cgdo = {5.932020000000001E-11/sw_func_tox_lv_ratio} cgbo = {0/sw_func_tox_lv_ratio}
+ ckappas = 0.6 cf = 1.2E-11 clc = 1E-7
+ cle = 0.6 dlc = -2.56E-9 dwc = 0
+ vfbcv = -0.1446893 noff = 4 voffcv = -0.1375
+ acde = 0.552 moin = 14.504 cgsl = {7.513892E-12/sw_func_tox_lv_ratio}
+ cgdl = {7.513892E-12/sw_func_tox_lv_ratio} ijthsrev = 0.1 ijthsfwd = 0.1
+ xjbvs = 1 bvs = 12.8 jss = 2.17E-5
+ jsws = 8.200000000000001E-10 cjs = {7.433E-04*sw_func_psd_nw_cj} mjs = 0.34629
+ mjsws = 0.26859 cjsws = {9.2435E-11*sw_func_psd_nw_cj} cjswgs = {2.4701E-10*sw_func_psd_nw_cj}
+ mjswgs = 0.70393 pbs = 0.6587 pbsws = 0.7418
+ pbswgs = 1.3925 xrcrg1 = 12 xrcrg2 = 1
+ rbpb = 50 rbpd = 50 rbps = 50
+ rbdb = 50 rbsb = 50 gbmin = 1E-12
+ tnom = 30 ute = -2.292033449469222 lute = 1.697840694396441E-5
+ wute = 1.388539590859364E-5 pute = -1.183950885889947E-10 kt1 = -0.438677016391383
+ lkt1 = -2.240114118306138E-7 wkt1 = 5.459594853740746E-8 pkt1 = 9.570625168036889E-13
+ kt1l = 0 kt2 = -0.046096682551354 lkt2 = 6.527681166444307E-8
+ wkt2 = 7.354565047893263E-8 pkt2 = -5.900949975307256E-13 ua1 = -4.901446257136616E-9
+ lua1 = 5.707166890506079E-14 wua1 = 4.820589450500103E-14 pua1 = -3.867809586787659E-19
+ ub1 = 4.303583952018314E-18 lub1 = -3.835995085217331E-23 wub1 = -3.436125864931392E-23
+ pub1 = 2.579844809775293E-28 uc1 = -8.842320167879033E-11 luc1 = 1.671084199133808E-15
+ wuc1 = 1.334140836749817E-15 puc1 = -1.07045056864789E-20 at = -4.630730766481792E5
+ lat = 3.715476091948199 wat = 1.389409387406994 pat = -1.114795400804776E-5
+ prt = 0 njs = 1.2556 xtis = 2
+ tpb = 1.9551E-3 tpbsw = 1.4242E-4 tpbswg = 0
+ tcj = 1.2407E-3 tcjsw = 0 tcjswg = 2E-12
+ tvoff = 0 tvfbsdoff = 0 saref = 3E-6
+ sbref = 3E-6 wlod = 0 ku0 = 4.5E-8
+ kvsat = 0.4 kvth0 = 2.65E-8 tku0 = 0
+ llodku0 = 0 wlodku0 = 1 llodvth = 0
+ wlodvth = 1 lku0 = 0 wku0 = 2.5E-7
+ pku0 = 0 lkvth0 = 0 wkvth0 = 2.5E-7
+ pkvth0 = 0 stk2 = 0 lodk2 = 1
+ steta0 = 0 lodeta0 = 1

.model phighvt_model.11 pmos
+ level = 54 lmin = 2E-6 lmax = 4E-6 wmin = 5E-6
+ wmax = 7E-6 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 4.23E-9
+ toxm = 4.23E-9 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 9.999999999999999E22 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {9.364E-9+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {-1.176E-8-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = -5.722E-9 dwb = -1.7864E-8 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = -1.132957133975123 lvth0 = 3.942346963175757E-8
+ wvth0 = 1.354075849398493E-7 pvth0 = -7.58509798024285E-14 k1 = 0.142984503762239
+ lk1 = 5.174534834031385E-7 wk1 = 1.541308769031606E-6 pk1 = -1.760654415458473E-12
+ k2 = 0.146679437452516 lk2 = -2.057690260441702E-7 wk2 = -6.064993416066668E-7
+ pk2 = 7.23317979983219E-13 k3 = -13.778 k3b = 2
+ w0 = 0 lpe0 = 0 lpeb = 0
+ vbm = -3 dvtp0 = 0 dvtp1 = 0
+ dvt0 = 4.05 dvt1 = 0.3 dvt2 = 0.03
+ dvt0w = -4.254 dvt1w = 1.1472E6 dvt2w = -8.96E-3
+ vfbsdoff = 0 u0 = 0.01938352761524 lu0 = -1.030904929347178E-8
+ wu0 = -3.358965328861184E-8 pu0 = 8.853896023498673E-15 ua = 9.921942718118987E-10
+ lua = -1.73337199594731E-15 wua = -5.150244343304943E-15 pua = -1.13813489172117E-21
+ ub = 3.725872679292201E-19 lub = 6.477203732166848E-25 wub = 1.52802365339835E-24
+ pub = 2.011833278753792E-30 uc = 7.102714358499673E-11 luc = -3.556953894138371E-16
+ wuc = -9.707123434556079E-16 puc = 2.415805928234238E-21 ud = 0
+ up = 0 lp = 1 eu = 1.67
+ vsat = 2.932006537212232E5 lvsat = -0.370331670408886 wvsat = -0.683767430907338
+ pvsat = 6.320536294899057E-7 a0 = 1.89451852078908 la0 = 5.183795805889164E-8
+ wa0 = -2.211924792239103E-7 pa0 = -2.382751365148178E-12 ags = 0.617032442091069
+ lags = 1.908867453667746E-7 wags = -8.901822445251887E-7 pags = 3.400790287840632E-12
+ b0 = 0 b1 = 0 keta = -0.087250574518802
+ lketa = 9.02240863894624E-8 wketa = 2.387936218399676E-7 pketa = -6.954705979858541E-13
+ a1 = 0 a2 = 0.8 rdsw = 531.92
+ rdswmin = 0 rdw = 0 rdwmin = 0
+ rsw = 0 rswmin = 0 prwb = -0.32348
+ prwg = 0.02 wr = 1 voff = -0.109847963959104
+ lvoff = -1.081631528476087E-7 wvoff = -5.672127748777806E-7 pvoff = 6.753504814686656E-13
+ voffl = 0 minv = 0 nfactor = 7.137640312840268
+ lnfactor = -7.049151852388439E-6 wnfactor = -2.934761488481259E-5 pnfactor = 3.586538125361819E-11
+ eta0 = 0.36076902740912 leta0 = -1.129679797161142E-6 weta0 = -1.398586894700282E-6
+ peta0 = 5.627242342564479E-12 etab = -0.31545216861552 letab = 9.87581709467917E-7
+ wetab = 1.222664014863769E-6 petab = -4.91941311708467E-12 dsub = 1.299735799480226
+ ldsub = -2.976341783924678E-6 wdsub = -3.684825225348463E-6 pdsub = 1.482596799069405E-11
+ cit = 1E-5 cdsc = 0 cdscb = 0
+ cdscd = 0 pclm = 0.272291943048333 lpclm = 1.45056167130617E-6
+ wpclm = 2.684505740238066E-6 ppclm = -1.080116253596267E-11 pdiblc1 = 0.39
+ pdiblc2 = 1.96039339360748E-3 lpdiblc2 = -3.32795753380188E-9 wpdiblc2 = -8.694279240561918E-9
+ ppdiblc2 = 1.657746168031636E-14 pdiblcb = 0.011424062641811 lpdiblcb = -2.62208359145415E-8
+ wpdiblcb = -7.970791950946565E-8 ppdiblcb = 1.612084133009103E-13 drout = 0.56
+ pscbe1 = 1.179482796167038E9 lpscbe1 = -765.2185455078293 wpscbe1 = -2.649272619362653E3
+ ppscbe1 = 5.342198805634534E-3 pscbe2 = 9.703400593916295E-9 lpscbe2 = -4.056067151511096E-15
+ wpscbe2 = -3.291311963480854E-15 ppscbe2 = 2.041328522579535E-20 pvag = 0
+ delta = 0.01 fprout = 0 pdits = 0
+ pditsl = 0 pditsd = 0 lambda = 0
+ vtl = 0 lc = 5E-9 xn = 3
+ alpha0 = 2.793180189910512E-3 lalpha0 = -1.123841595535674E-8 walpha0 = -1.949994995264974E-8
+ palpha0 = 7.845843863348529E-14 alpha1 = -1.519925879360001E-10 lalpha1 = 1.013897217412255E-15
+ walpha1 = 1.759228798365135E-15 palpha1 = -7.078292254798087E-21 beta0 = 68.04964503300299
+ lbeta0 = -2.589428905393242E-4 wbeta0 = -4.519113846103392E-4 pbeta0 = 1.86389379955358E-9
+ aigbacc = 0.43 bigbacc = 0.054 cigbacc = 0.075
+ nigbacc = 1 aigbinv = 0.35 bigbinv = 0.03
+ cigbinv = 6E-3 eigbinv = 1.1 nigbinv = 3
+ aigc = 0.43 bigc = 0.054 cigc = 0.075
+ aigsd = 0.43 bigsd = 0.054 cigsd = 0.075
+ dlcig = 0 nigc = 1 poxedge = 1
+ pigcd = 1 ntox = 1 toxref = 4.23E-9
+ agidl = -1.836148507089743E-8 lagidl = 3.739446488807231E-14 wagidl = 1.294841321101976E-13
+ pagidl = -2.62199435903274E-19 bgidl = -3.303865438217136E9 lbgidl = 7.02472299531611E3
+ wbgidl = 3.004645527559302E4 pbgidl = -0.049041501954956 cgidl = 300
+ egidl = -0.951128598301789 legidl = 2.126979741235637E-6 wegidl = 7.33821465172353E-6
+ pegidl = -1.48490241120556E-11 noia = 1.2E41 noib = 2E25
+ noic = 0 em = 4.1E7 af = 1
+ ef = 0.88 kf = 0 lintnoi = -6E-8
+ tnoia = 1.5 tnoib = 3.5 ntnoi = 1
+ rnoia = 0.577 rnoib = 0.37 xpart = 0
+ cgso = {5.932020000000001E-11/sw_func_tox_lv_ratio} cgdo = {5.932020000000001E-11/sw_func_tox_lv_ratio} cgbo = {0/sw_func_tox_lv_ratio}
+ ckappas = 0.6 cf = 1.2E-11 clc = 1E-7
+ cle = 0.6 dlc = -2.56E-9 dwc = 0
+ vfbcv = -0.1446893 noff = 4 voffcv = -0.1375
+ acde = 0.552 moin = 14.504 cgsl = {7.513892E-12/sw_func_tox_lv_ratio}
+ cgdl = {7.513892E-12/sw_func_tox_lv_ratio} ijthsrev = 0.1 ijthsfwd = 0.1
+ xjbvs = 1 bvs = 12.8 jss = 2.17E-5
+ jsws = 8.200000000000001E-10 cjs = {7.433E-04*sw_func_psd_nw_cj} mjs = 0.34629
+ mjsws = 0.26859 cjsws = {9.2435E-11*sw_func_psd_nw_cj} cjswgs = {2.4701E-10*sw_func_psd_nw_cj}
+ mjswgs = 0.70393 pbs = 0.6587 pbsws = 0.7418
+ pbswgs = 1.3925 xrcrg1 = 12 xrcrg2 = 1
+ rbpb = 50 rbpd = 50 rbps = 50
+ rbdb = 50 rbsb = 50 gbmin = 1E-12
+ tnom = 30 ute = 4.296448953374693 lute = -9.53048377352614E-6
+ wute = -3.300664421982667E-5 pute = 7.027597270850702E-11 kt1 = -0.588402303620551
+ lkt1 = 3.784112758416892E-7 wkt1 = 7.951393272591422E-7 pkt1 = -2.022528578350785E-12
+ kt1l = 0 kt2 = -0.029528643749617 lkt2 = -1.385023815121792E-9
+ wkt2 = -5.187073765662651E-8 pkt2 = -8.547965153954073E-14 ua1 = 1.782893088620175E-8
+ lua1 = -3.438445813870399E-14 wua1 = -1.0346574937129E-13 pua1 = 2.234729338903684E-19
+ ub1 = -1.144795964250754E-17 lub1 = 2.501669983127332E-23 wub1 = 7.082446911122874E-23
+ pub1 = -1.652323983815693E-28 uc1 = 1.050703613276522E-9 luc1 = -2.912215323375188E-15
+ wuc1 = -4.90146736349043E-15 puc1 = 1.438458861935174E-20 at = 7.388026945837544E5
+ lat = -1.120295111118911 wat = -2.112983624988177 pat = 2.943994325184456E-6
+ prt = 0 njs = 1.2556 xtis = 2
+ tpb = 1.9551E-3 tpbsw = 1.4242E-4 tpbswg = 0
+ tcj = 1.2407E-3 tcjsw = 0 tcjswg = 2E-12
+ tvoff = 0 tvfbsdoff = 0 saref = 3E-6
+ sbref = 3E-6 wlod = 0 ku0 = 4.5E-8
+ kvsat = 0.4 kvth0 = 2.65E-8 tku0 = 0
+ llodku0 = 0 wlodku0 = 1 llodvth = 0
+ wlodvth = 1 lku0 = 0 wku0 = 2.5E-7
+ pku0 = 0 lkvth0 = 0 wkvth0 = 2.5E-7
+ pkvth0 = 0 stk2 = 0 lodk2 = 1
+ steta0 = 0 lodeta0 = 1

.model phighvt_model.12 pmos
+ level = 54 lmin = 1E-6 lmax = 2E-6 wmin = 5E-6
+ wmax = 7E-6 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 4.23E-9
+ toxm = 4.23E-9 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 9.999999999999999E22 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {9.364E-9+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {-1.176E-8-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = -5.722E-9 dwb = -1.7864E-8 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = -1.146553362234986 lvth0 = 6.693570944015578E-8
+ wvth0 = 2.267587057383265E-7 pvth0 = -2.607017997605632E-13 k1 = 0.343329859335146
+ lk1 = 1.120506494942503E-7 wk1 = 1.416868582927932E-6 pk1 = -1.508847210073965E-12
+ k2 = 0.060368423255552 lk2 = -3.111696259632864E-8 wk2 = -4.79475153296175E-7
+ pk2 = 4.662819944531725E-13 k3 = -13.778 k3b = 2
+ w0 = 0 lpe0 = 0 lpeb = 0
+ vbm = -3 dvtp0 = 0 dvtp1 = 0
+ dvt0 = 4.05 dvt1 = 0.3 dvt2 = 0.03
+ dvt0w = -4.254 dvt1w = 1.1472E6 dvt2w = -8.96E-3
+ vfbsdoff = 0 u0 = 0.018388893136669 lu0 = -8.296386533393471E-9
+ wu0 = -5.73796598486667E-8 pu0 = 5.699345009790088E-14 ua = 1.002142238646745E-9
+ lua = -1.753501905796959E-15 wua = -1.197800772656341E-14 pua = 1.267798086957001E-20
+ ub = 2.8922459203206E-19 lub = 8.164064151481064E-25 wub = 5.776618352224E-24
+ pub = -6.585283066213888E-30 uc = -1.279682227409016E-10 luc = 4.697571425394468E-17
+ wuc = 3.221670275954014E-16 puc = -2.003613366748999E-22 ud = 0
+ up = 0 lp = 1 eu = 1.67
+ vsat = 9.123788455499537E4 lvsat = 0.03834403225436 wvsat = -0.466098237497293
+ pvsat = 1.915956632408128E-7 a0 = 0.704598172126722 la0 = 2.459665581984146E-6
+ wa0 = 7.2258321063797E-6 pa0 = -1.74519545546088E-11 ags = -0.534717359631118
+ lags = 2.521475504147655E-6 wags = 8.389232316470883E-6 pags = -1.537629066462614E-11
+ b0 = 0 b1 = 0 keta = 0.028793478633901
+ lketa = -1.445933760460949E-7 wketa = -7.163754193400901E-7 pketa = 1.237333060222816E-12
+ a1 = 0 a2 = 0.8 rdsw = 531.92
+ rdswmin = 0 rdw = 0 rdwmin = 0
+ rsw = 0 rswmin = 0 prwb = -0.32348
+ prwg = 0.02 wr = 1 voff = -0.12244647675584
+ lvoff = -8.266981023315802E-8 wvoff = -4.613655431939578E-7 pvoff = 4.611664912118166E-13
+ voffl = 0 minv = 0 nfactor = 6.17445676774314
+ lnfactor = -5.100130685213499E-6 wnfactor = -2.581386354078717E-5 pnfactor = 2.871476473395587E-11
+ eta0 = -0.624049819054026 leta0 = 8.631208350339629E-7 weta0 = 2.793283237817287E-6
+ peta0 = -2.855090707987473E-12 etab = -0.421273590909305 letab = 1.201713473907836E-6
+ wetab = 2.941107624313303E-6 petab = -8.396718129677993E-12 dsub = -1.74362717546396
+ ldsub = 3.18196406313438E-6 wdsub = 9.979297232911128E-6 pdsub = -1.28236570860434E-11
+ cit = 1E-5 cdsc = 0 cdscb = 0
+ cdscd = 0 pclm = 0.962044522764335 lpclm = 5.483353119924648E-8
+ wpclm = -3.271031405718408E-6 ppclm = 1.249985989623181E-12 pdiblc1 = 0.536396434431536
+ lpdiblc1 = -2.962361130009008E-7 wpdiblc1 = -6.972946565473529E-7 ppdiblc1 = 1.4109896834167E-12
+ pdiblc2 = 1.988241060307262E-4 lpdiblc2 = 2.366131509954311E-10 wpdiblc2 = -1.015586248545487E-9
+ ppdiblc2 = 1.039472837111277E-15 pdiblcb = -0.062046077268656 lpdiblcb = 1.224474615970882E-7
+ wpdiblcb = 4.209850679957316E-7 ppdiblcb = -8.519538607756064E-13 drout = -0.110414672003951
+ ldrout = 1.356597497093435E-6 wdrout = 2.612387484578341E-6 pdrout = -5.286218322793964E-12
+ pscbe1 = 7.9946973E8 pscbe2 = 6.529375979152383E-9 lpscbe2 = 2.366635136955977E-15
+ wpscbe2 = 1.187688649718058E-14 ppscbe2 = -1.027986772332229E-20 pvag = 0
+ delta = 0.01 fprout = 0 pdits = 0
+ pditsl = 0 pditsd = 0 lambda = 0
+ vtl = 0 lc = 5E-9 xn = 3
+ alpha0 = -5.550299118422882E-3 lalpha0 = 5.644781294642048E-9 walpha0 = 3.874814852519756E-8
+ palpha0 = -3.940775359840829E-14 alpha1 = 3.490636E-10 walpha1 = -1.7387807368992E-15
+ beta0 = -81.13928659192514 lbeta0 = 4.294389638235034E-5 wbeta0 = 6.065013584500198E-4
+ pbeta0 = -2.778255542839178E-10 aigbacc = 0.43 bigbacc = 0.054
+ cigbacc = 0.075 nigbacc = 1 aigbinv = 0.35
+ bigbinv = 0.03 cigbinv = 6E-3 eigbinv = 1.1
+ nigbinv = 3 aigc = 0.43 bigc = 0.054
+ cigc = 0.075 aigsd = 0.43 bigsd = 0.054
+ cigsd = 0.075 dlcig = 0 nigc = 1
+ poxedge = 1 pigcd = 1 ntox = 1
+ toxref = 4.23E-9 agidl = 1.372806174099593E-10 lagidl = -3.815745753144158E-17
+ wagidl = -1.85704895646943E-16 pagidl = 1.900726747925591E-22 bgidl = -1.17651291172094E8
+ lbgidl = 577.3549444875264 wbgidl = 6.89846042087413E3 pbgidl = -2.201071406535717E-3
+ cgidl = 300 egidl = 0.1 noia = 1.2E41
+ noib = 2E25 noic = 0 em = 4.1E7
+ af = 1 ef = 0.88 kf = 0
+ lintnoi = -6E-8 tnoia = 1.5 tnoib = 3.5
+ ntnoi = 1 rnoia = 0.577 rnoib = 0.37
+ xpart = 0 cgso = {5.932020000000001E-11/sw_func_tox_lv_ratio} cgdo = {5.932020000000001E-11/sw_func_tox_lv_ratio}
+ cgbo = {0/sw_func_tox_lv_ratio} ckappas = 0.6 cf = 1.2E-11
+ clc = 1E-7 cle = 0.6 dlc = -2.56E-9
+ dwc = 0 vfbcv = -0.1446893 noff = 4
+ voffcv = -0.1375 acde = 0.552 moin = 14.504
+ cgsl = {7.513892E-12/sw_func_tox_lv_ratio} cgdl = {7.513892E-12/sw_func_tox_lv_ratio} ijthsrev = 0.1
+ ijthsfwd = 0.1 xjbvs = 1 bvs = 12.8
+ jss = 2.17E-5 jsws = 8.200000000000001E-10 cjs = {7.433E-04*sw_func_psd_nw_cj}
+ mjs = 0.34629 mjsws = 0.26859 cjsws = {9.2435E-11*sw_func_psd_nw_cj}
+ cjswgs = {2.4701E-10*sw_func_psd_nw_cj} mjswgs = 0.70393 pbs = 0.6587
+ pbsws = 0.7418 pbswgs = 1.3925 xrcrg1 = 12
+ xrcrg2 = 1 rbpb = 50 rbpd = 50
+ rbps = 50 rbdb = 50 rbsb = 50
+ gbmin = 1E-12 tnom = 30 ute = 0.547694456095267
+ lute = -1.944804073191279E-6 wute = 3.902303394421914E-6 pute = -4.410020967877276E-12
+ kt1 = -0.353992558099684 lkt1 = -9.592153241469436E-8 wkt1 = -2.480014595800781E-7
+ pkt1 = 8.828766663411361E-14 kt1l = 0 kt2 = -0.01126756896176
+ lkt2 = -3.833667386984657E-8 wkt2 = -2.014245981073796E-7 pkt2 = 2.171455761597671E-13
+ ua1 = 3.005299628336953E-9 lua1 = -4.388543815789414E-15 wua1 = 9.552943512643646E-15
+ pua1 = -5.22265153412888E-21 ub1 = -5.867946439504858E-20 lub1 = 1.970263605259153E-24
+ wub1 = -1.404345509933589E-23 pub1 = 6.499543616992422E-30 uc1 = -6.996263011071186E-10
+ luc1 = 6.29612264978395E-16 wuc1 = 3.864418818298844E-15 puc1 = -3.353357387222486E-21
+ at = 1.295071729805303E5 lat = 0.112626562755645 wat = -0.666194307713501
+ pat = 1.638720589280301E-8 prt = 0 njs = 1.2556
+ xtis = 2 tpb = 1.9551E-3 tpbsw = 1.4242E-4
+ tpbswg = 0 tcj = 1.2407E-3 tcjsw = 0
+ tcjswg = 2E-12 tvoff = 0 tvfbsdoff = 0
+ saref = 3E-6 sbref = 3E-6 wlod = 0
+ ku0 = 4.5E-8 kvsat = 0.4 kvth0 = 2.65E-8
+ tku0 = 0 llodku0 = 0 wlodku0 = 1
+ llodvth = 0 wlodvth = 1 lku0 = 0
+ wku0 = 2.5E-7 pku0 = 0 lkvth0 = 0
+ wkvth0 = 2.5E-7 pkvth0 = 0 stk2 = 0
+ lodk2 = 1 steta0 = 0 lodeta0 = 1

.model phighvt_model.13 pmos
+ level = 54 lmin = 5E-7 lmax = 1E-6 wmin = 5E-6
+ wmax = 7E-6 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 4.23E-9
+ toxm = 4.23E-9 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 9.999999999999999E22 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {9.364E-9+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {-1.176E-8-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = -5.722E-9 dwb = -1.7864E-8 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = -1.070756495030402 lvth0 = -1.064390008108057E-8
+ wvth0 = -2.310222788989885E-7 pvth0 = 2.078461936354215E-13 k1 = 0.435301124941151
+ lk1 = 1.79162197211924E-8 wk1 = -1.895122268194113E-7 pk1 = 1.353156763186348E-13
+ k2 = 0.044309254926654 lk2 = -1.468008262833541E-8 wk2 = -4.009275317217974E-8
+ pk2 = 1.656532027826102E-14 k3 = -13.778 k3b = 2
+ w0 = 0 lpe0 = 0 lpeb = 0
+ vbm = -3 dvtp0 = 0 dvtp1 = 0
+ dvt0 = 4.05 dvt1 = 0.3 dvt2 = 0.03
+ dvt0w = -4.254 dvt1w = 1.1472E6 dvt2w = -8.96E-3
+ vfbsdoff = 0 u0 = 0.010147423756238 lu0 = 1.389222068651935E-10
+ wu0 = 1.568771443226841E-8 pu0 = -1.779246882612182E-14 ua = -6.8378595726444E-10
+ lua = -2.792067871794308E-17 wua = 3.977202204860707E-15 pua = -3.652495599441205E-21
+ ub = 1.060784935026221E-18 lub = 2.66989728867226E-26 wub = -2.519209647726477E-24
+ pub = 1.905662808295423E-30 uc = -1.416036311715854E-10 luc = 6.09318274909182E-17
+ wuc = 1.832844893417354E-16 puc = -5.821228112150779E-23 ud = 0
+ up = 0 lp = 1 eu = 1.67
+ vsat = 1.800767740652203E5 lvsat = -0.052584347937146 wvsat = -0.77401532583204
+ pvsat = 5.067549614931922E-7 a0 = 5.709227320964977 la0 = -2.662672444434784E-6
+ wa0 = -2.348040177228553E-5 pa0 = 1.397648994488264E-11 ags = 3.401465835451707
+ lags = -1.507286719683517E-6 wags = -1.65970869270733E-5 pags = 1.01977068075262E-11
+ b0 = 0 b1 = 0 keta = -0.20190732069733
+ lketa = 9.153350608540654E-8 wketa = 1.035234285103897E-6 pketa = -5.554745044696932E-13
+ a1 = 0 a2 = 0.150625341882111 la2 = 6.646479500768218E-7
+ wa2 = 3.071526911251993E-6 pa2 = -3.143769224204639E-12 rdsw = 531.92
+ rdswmin = 0 rdw = 0 rdwmin = 0
+ rsw = 0 rswmin = 0 prwb = -0.32348
+ prwg = 0.02 wr = 1 voff = -0.292038930652971
+ lvoff = 9.091145817963288E-8 wvoff = 5.136576603086495E-7 pvoff = -5.367892580371718E-13
+ voffl = 0 minv = 0 nfactor = -4.80746467992791
+ lnfactor = 6.140085554906772E-6 wnfactor = 3.472481369420692E-5 pnfactor = -3.324778218960527E-11
+ eta0 = 0.540016491075685 leta0 = -3.283243147099987E-7 weta0 = -7.328047010929604E-7
+ peta0 = 7.539308192459435E-13 etab = 1.544391920644272 letab = -8.101844904774806E-7
+ wetab = -1.078880134462008E-5 petab = 5.656118298204702E-12 dsub = 1.747613553007017
+ ldsub = -3.913906472702334E-7 wdsub = -5.219293564428404E-6 pdsub = 2.732404566849558E-12
+ cit = 1E-5 cdsc = 0 cdscb = 0
+ cdscd = 0 pclm = 0.474665005454713 lpclm = 5.536762147559903E-7
+ wpclm = 5.050522221713854E-7 ppclm = -2.614911125194581E-12 pdiblc1 = 1.335071146741042
+ lpdiblc1 = -1.113695654543927E-6 wpdiblc1 = -4.804314372447336E-6 ppdiblc1 = 5.61460650303465E-12
+ pdiblc2 = 2.229783483387561E-3 lpdiblc2 = -1.842114390916836E-9 wpdiblc2 = -1.509865276980028E-8
+ ppdiblc2 = 1.545377308294598E-14 pdiblcb = 0.144060121182146 lpdiblcb = -8.850635464127708E-8
+ wpdiblcb = -8.421344479612309E-7 ppdiblcb = 4.408742261966636E-13 drout = 0.845234810612308
+ ldrout = 3.784711386460419E-7 wdrout = -7.297870108350228E-7 pdrout = -1.865435883248478E-12
+ pscbe1 = 9.499741652986158E8 lpscbe1 = -153.50155766643925 wpscbe1 = -747.0621103253667
+ ppscbe1 = 7.646330111602193E-4 pscbe2 = 8.944163671910632E-9 lpscbe2 = -1.049483623359464E-16
+ wpscbe2 = 8.893600509951148E-16 ppscbe2 = 9.660853448774623E-22 pvag = 0
+ delta = 0.01 fprout = 0 pdits = 0
+ pditsl = 0 pditsd = 0 lambda = 0
+ vtl = 0 lc = 5E-9 xn = 3
+ alpha0 = -7.212182279628058E-5 lalpha0 = 3.775726902230881E-11 walpha0 = 5.035027602038354E-10
+ palpha0 = -2.635937650219119E-16 alpha1 = 6.098431517439999E-10 lalpha1 = -2.669130868010188E-16
+ walpha1 = -3.559353719662139E-15 palpha1 = 1.863392859317523E-21 beta0 = -89.49517053003437
+ lbeta0 = 5.149631071068392E-5 wbeta0 = 6.844222939640521E-4 pbeta0 = -3.5757919020124E-10
+ aigbacc = 0.43 bigbacc = 0.054 cigbacc = 0.075
+ nigbacc = 1 aigbinv = 0.35 bigbinv = 0.03
+ cigbinv = 6E-3 eigbinv = 1.1 nigbinv = 3
+ aigc = 0.43 bigc = 0.054 cigc = 0.075
+ aigsd = 0.43 bigsd = 0.054 cigsd = 0.075
+ dlcig = 0 nigc = 1 poxedge = 1
+ pigcd = 1 ntox = 1 toxref = 4.23E-9
+ agidl = 1E-10 bgidl = -3.220042722822843E8 lbgidl = 786.5143077134283
+ wbgidl = 9.801451347878769E3 pbgidl = -5.172340680143504E-3 cgidl = 300
+ egidl = 0.1 noia = 1.2E41 noib = 2E25
+ noic = 0 em = 4.1E7 af = 1
+ ef = 0.88 kf = 0 lintnoi = -6E-8
+ tnoia = 1.5 tnoib = 3.5 ntnoi = 1
+ rnoia = 0.577 rnoib = 0.37 xpart = 0
+ cgso = {5.932020000000001E-11/sw_func_tox_lv_ratio} cgdo = {5.932020000000001E-11/sw_func_tox_lv_ratio} cgbo = {0/sw_func_tox_lv_ratio}
+ ckappas = 0.6 cf = 1.2E-11 clc = 1E-7
+ cle = 0.6 dlc = -2.56E-9 dwc = 0
+ vfbcv = -0.1446893 noff = 4 voffcv = -0.1375
+ acde = 0.552 moin = 14.504 cgsl = {7.513892E-12/sw_func_tox_lv_ratio}
+ cgdl = {7.513892E-12/sw_func_tox_lv_ratio} ijthsrev = 0.1 ijthsfwd = 0.1
+ xjbvs = 1 bvs = 12.8 jss = 2.17E-5
+ jsws = 8.200000000000001E-10 cjs = {7.433E-04*sw_func_psd_nw_cj} mjs = 0.34629
+ mjsws = 0.26859 cjsws = {9.2435E-11*sw_func_psd_nw_cj} cjswgs = {2.4701E-10*sw_func_psd_nw_cj}
+ mjswgs = 0.70393 pbs = 0.6587 pbsws = 0.7418
+ pbswgs = 1.3925 xrcrg1 = 12 xrcrg2 = 1
+ rbpb = 50 rbpd = 50 rbps = 50
+ rbdb = 50 rbsb = 50 gbmin = 1E-12
+ tnom = 30 ute = -2.653281286977302 lute = 1.331458619358357E-6
+ wute = -8.318707952371187E-7 pute = 4.355009987225364E-13 kt1 = -0.405500572067165
+ lkt1 = -4.320204995869872E-8 wkt1 = -3.138867931185881E-7 pkt1 = 1.557226232174494E-13
+ kt1l = 0 kt2 = -0.069612872533422 lkt2 = 2.138091124182081E-8
+ wkt2 = 5.042262617049748E-8 pkt2 = -4.062509483312558E-14 ua1 = -5.460209246226802E-9
+ lua1 = 4.276073827504079E-15 wua1 = 1.014221930109088E-14 pua1 = -5.825787089120392E-21
+ ub1 = 6.418331373203003E-18 lub1 = -4.659086527239203E-24 wub1 = -1.865042042708382E-23
+ pub1 = 1.121486476924898E-29 uc1 = 6.646302349651712E-11 luc1 = -1.544954805399182E-16
+ wuc1 = 9.60368896034277E-16 puc1 = -3.81004210786257E-22 at = 4.762483033545739E5
+ lat = -0.242269919004796 wat = -1.524824800810664 pat = 8.952126881876115E-7
+ prt = 0 njs = 1.2556 xtis = 2
+ tpb = 1.9551E-3 tpbsw = 1.4242E-4 tpbswg = 0
+ tcj = 1.2407E-3 tcjsw = 0 tcjswg = 2E-12
+ tvoff = 0 tvfbsdoff = 0 saref = 2.75E-6
+ sbref = 2.74E-6 wlod = 0 ku0 = 4.5E-8
+ kvsat = 0.4 kvth0 = 2.65E-8 tku0 = 0
+ llodku0 = 0 wlodku0 = 1 llodvth = 0
+ wlodvth = 1 lku0 = 0 wku0 = 2.5E-7
+ pku0 = 0 lkvth0 = 0 wkvth0 = 2.5E-7
+ pkvth0 = 0 stk2 = 0 lodk2 = 1
+ steta0 = 0 lodeta0 = 1

.model phighvt_model.14 pmos
+ level = 54 lmin = 2.5E-7 lmax = 5E-7 wmin = 5E-6
+ wmax = 7E-6 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 4.23E-9
+ toxm = 4.23E-9 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 9.999999999999999E22 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {9.364E-9+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {-1.176E-8-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = -5.722E-9 dwb = -1.7864E-8 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = -1.112364947487036 lvth0 = 1.11389569490168E-8
+ wvth0 = 2.638597186502858E-7 pvth0 = -5.123442972157464E-14 k1 = 0.201650054649689
+ lk1 = 1.402372280401785E-7 wk1 = -1.063149960990127E-7 pk1 = 9.176026209189169E-14
+ k2 = 0.104108427891092 lk2 = -4.598614565867784E-8 wk2 = 8.58020668609849E-8
+ pk2 = -4.934313590550132E-14 k3 = -13.778 k3b = 2
+ w0 = 0 lpe0 = 0 lpeb = 0
+ vbm = -3 dvtp0 = 0 dvtp1 = 0
+ dvt0 = 4.05 dvt1 = 0.3 dvt2 = 0.03
+ dvt0w = -4.254 dvt1w = 1.1472E6 dvt2w = -8.96E-3
+ vfbsdoff = 0 u0 = 0.016624234646526 lu0 = -3.251817830418588E-9
+ wu0 = -3.886566650591568E-8 pu0 = 1.076731716263632E-14 ua = 6.662618482508327E-10
+ lua = -7.346977058612986E-16 wua = -7.368621654057315E-15 pua = 2.287270107179558E-21
+ ub = 3.314638056780336E-19 lub = 4.085131705230856E-25 wub = 3.285899257005749E-24
+ pub = -1.133427805509991E-30 uc = -8.98050151379466E-11 luc = 3.381421602498762E-17
+ wuc = 4.091354543185826E-16 puc = -1.764497783061868E-22 ud = 0
+ up = 0 lp = 1 eu = 1.67
+ vsat = 8.410823663606925E4 lvsat = -2.342899222236581E-3 wvsat = 0.351817355507319
+ pvsat = -8.264096384158857E-8 a0 = 0.346533311530829 la0 = 1.448051233841804E-7
+ wa0 = 7.454072673506576E-6 pa0 = -2.218326116978446E-12 ags = -2.364577166002175
+ lags = 1.511352112437619E-6 wags = 1.256411690250589E-5 pags = -5.0687666213351E-12
+ b0 = 0 b1 = 0 keta = 3.954702331472652E-3
+ lketa = -1.623938021063208E-8 wketa = 1.910090589709981E-7 pketa = -1.13505714084598E-13
+ a1 = 0 a2 = 2.098749316235778 la2 = -3.552339129768099E-7
+ wa2 = -6.143053822503984E-6 pa2 = 1.680248081531289E-12 rdsw = 531.92
+ rdswmin = 0 rdw = 0 rdwmin = 0
+ rsw = 0 rswmin = 0 prwb = -0.32348
+ prwg = 0.02 wr = 1 voff = -0.021023265217025
+ lvoff = -5.097066298939347E-8 wvoff = -9.295573593398337E-7 pvoff = 2.18762669049202E-13
+ voffl = 0 minv = 0 nfactor = 11.433594687342344
+ lnfactor = -2.36243384504655E-6 wnfactor = -5.357878463859777E-5 pnfactor = 1.298091760958464E-11
+ eta0 = -0.718558725208225 leta0 = 3.305649825189536E-7 weta0 = 1.481171608519028E-6
+ peta0 = -4.051300583621244E-13 etab = -5.973928727164705E-3 letab = 1.46303898545409E-9
+ wetab = 3.186007307679059E-8 petab = -8.714367187963762E-15 dsub = 1.450662922633179
+ ldsub = -2.359310532569218E-7 wdsub = -7.288921885309258E-7 pdsub = 3.815896385397103E-13
+ cit = 1E-5 cdsc = 0 cdscb = 0
+ cdscd = 0 pclm = 2.188538802492949 lpclm = -3.435709954694669E-7
+ wpclm = -7.796048968549642E-6 ppclm = 1.730881370171691E-12 pdiblc1 = -2.214995844492069
+ lpdiblc1 = 7.448354167064313E-7 wpdiblc1 = 1.341626180508516E-5 ppdiblc1 = -3.924229537427162E-12
+ pdiblc2 = -0.011803611726047 lpdiblc2 = 5.504648669126206E-9 wpdiblc2 = 2.905856683503168E-8
+ ppdiblc2 = -7.663414524575645E-15 pdiblcb = -0.025 drout = 2.347480819751035
+ ldrout = -4.079846920582645E-7 wdrout = -6.746513368502991E-6 pdrout = 1.284440699517856E-12
+ pscbe1 = 5.000516694027684E8 lpscbe1 = 82.04186738495478 wpscbe1 = 1.494124220650733E3
+ ppscbe1 = -4.086728568323885E-4 pscbe2 = 1.721592081273083E-8 lpscbe2 = -4.435378660698136E-15
+ wpscbe2 = 5.726732475097699E-15 ppscbe2 = -1.566375866588723E-21 pvag = 0
+ delta = 0.01 fprout = 0 pdits = 0
+ pditsl = 0 pditsd = 0 lambda = 0
+ vtl = 0 lc = 5E-9 xn = 3
+ alpha0 = -5.9785822459679E-8 lalpha0 = 3.135142577409115E-14 walpha0 = 2.983075706153702E-13
+ palpha0 = -1.561699793685586E-19 alpha1 = 4.819035034879999E-10 lalpha1 = -1.999341221460377E-16
+ walpha1 = -1.902365228626677E-15 palpha1 = 9.959262444906377E-22 beta0 = -20.978583903706497
+ lbeta0 = 1.562650728006875E-5 wbeta0 = 1.518878596266096E-4 pbeta0 = -7.878676313690216E-11
+ aigbacc = 0.43 bigbacc = 0.054 cigbacc = 0.075
+ nigbacc = 1 aigbinv = 0.35 bigbinv = 0.03
+ cigbinv = 6E-3 eigbinv = 1.1 nigbinv = 3
+ aigc = 0.43 bigc = 0.054 cigc = 0.075
+ aigsd = 0.43 bigsd = 0.054 cigsd = 0.075
+ dlcig = 0 nigc = 1 poxedge = 1
+ pigcd = 1 ntox = 1 toxref = 4.23E-9
+ agidl = 1E-10 bgidl = 9.928906596336955E8 lbgidl = 98.14051295677457
+ wbgidl = 671.2896635880518 pbgidl = -3.925184351836281E-4 cgidl = 300
+ egidl = 0.1 noia = 1.2E41 noib = 2E25
+ noic = 0 em = 4.1E7 af = 1
+ ef = 0.88 kf = 0 lintnoi = -6E-8
+ tnoia = 1.5 tnoib = 3.5 ntnoi = 1
+ rnoia = 0.577 rnoib = 0.37 xpart = 0
+ cgso = {5.932020000000001E-11/sw_func_tox_lv_ratio} cgdo = {5.932020000000001E-11/sw_func_tox_lv_ratio} cgbo = {0/sw_func_tox_lv_ratio}
+ ckappas = 0.6 cf = 1.2E-11 clc = 1E-7
+ cle = 0.6 dlc = -2.56E-9 dwc = 0
+ vfbcv = -0.1446893 noff = 4 voffcv = -0.1375
+ acde = 0.552 moin = 14.504 cgsl = {7.513892E-12/sw_func_tox_lv_ratio}
+ cgdl = {7.513892E-12/sw_func_tox_lv_ratio} ijthsrev = 0.1 ijthsfwd = 0.1
+ xjbvs = 1 bvs = 12.8 jss = 2.17E-5
+ jsws = 8.200000000000001E-10 cjs = {7.433E-04*sw_func_psd_nw_cj} mjs = 0.34629
+ mjsws = 0.26859 cjsws = {9.2435E-11*sw_func_psd_nw_cj} cjswgs = {2.4701E-10*sw_func_psd_nw_cj}
+ mjswgs = 0.70393 pbs = 0.6587 pbsws = 0.7418
+ pbswgs = 1.3925 xrcrg1 = 12 xrcrg2 = 1
+ rbpb = 50 rbpd = 50 rbps = 50
+ rbdb = 50 rbsb = 50 gbmin = 1E-12
+ tnom = 30 ute = -0.11297083419776 lute = 1.555291119211311E-9
+ wute = -4.375440025841357E-7 pute = 2.290630362328467E-13 kt1 = -0.425251065137649
+ lkt1 = -3.286227182643905E-8 wkt1 = -4.049357165514104E-7 pkt1 = 2.033885556130005E-13
+ kt1l = 0 kt2 = -0.023202834500706 lkt2 = -2.915671869066648E-9
+ wkt2 = -2.247145986094128E-8 pkt2 = -2.463582913946768E-15 ua1 = 4.427681481291919E-9
+ lua1 = -9.004347261665214E-16 wua1 = -2.579239405806088E-15 pua1 = 8.341509731143098E-22
+ ub1 = -4.781699272733067E-18 lub1 = 1.204353516521247E-24 wub1 = 8.587119984942831E-24
+ pub1 = -3.044532387255208E-30 uc1 = -3.387452461729892E-10 luc1 = 5.763915279746179E-17
+ wuc1 = 7.557584604882635E-17 puc1 = 8.220264674212598E-23 at = -4.305382274874838E4
+ lat = 0.029595130052815 wat = 0.539439247969623 pat = -1.854708266298443E-7
+ prt = 0 njs = 1.2556 xtis = 2
+ tpb = 1.9551E-3 tpbsw = 1.4242E-4 tpbswg = 0
+ tcj = 1.2407E-3 tcjsw = 0 tcjswg = 2E-12
+ tvoff = 0 tvfbsdoff = 0 saref = 1.75E-6
+ sbref = 1.74E-6 wlod = 0 ku0 = 4.5E-8
+ kvsat = 0.4 kvth0 = 2.65E-8 tku0 = 0
+ llodku0 = 0 wlodku0 = 1 llodvth = 0
+ wlodvth = 1 lku0 = 0 wku0 = 2.5E-7
+ pku0 = 0 lkvth0 = 0 wkvth0 = 2.5E-7
+ pkvth0 = 0 stk2 = 0 lodk2 = 1
+ steta0 = 0 lodeta0 = 1

.model phighvt_model.15 pmos
+ level = 54 lmin = 1.8E-7 lmax = 2.5E-7 wmin = 5E-6
+ wmax = 7E-6 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 4.23E-9
+ toxm = 4.23E-9 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 9.999999999999999E22 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {9.364E-9+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {-1.176E-8-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = -5.722E-9 dwb = -1.7864E-8 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = -1.071553779454965 lvth0 = -2.371373111523413E-11
+ wvth0 = 5.422917827619508E-7 pvth0 = -1.273911678973973E-13 k1 = -0.717901943764421
+ lk1 = 3.917530906464059E-7 wk1 = 5.419422020076108E-6 pk1 = -1.419639326572327E-12
+ k2 = 0.454717842960246 lk2 = -1.418848328683929E-7 wk2 = -1.829933284557793E-6
+ pk2 = 4.746487974145628E-13 k3 = -13.778 k3b = 2
+ w0 = 0 lpe0 = 0 lpeb = 0
+ vbm = -3 dvtp0 = 0 dvtp1 = 0
+ dvt0 = 4.05 dvt1 = 0.3 dvt2 = 0.03
+ dvt0w = -4.254 dvt1w = 1.1472E6 dvt2w = -8.96E-3
+ vfbsdoff = 0 u0 = 0.025294696068799 lu0 = -5.623362438638718E-9
+ wu0 = -1.140700215924584E-7 pu0 = 3.133721236590748E-14 ua = 3.87696302797749E-9
+ lua = -1.612888692540134E-15 wua = -3.190874690658725E-14 pua = 8.999485166251544E-21
+ ub = -2.324599821110689E-18 lub = 1.134999693722337E-24 wub = 2.239333083103938E-23
+ pub = -6.35969248963967E-30 uc = 6.986948200804822E-11 luc = -9.859952434384879E-18
+ wuc = -2.651716403380722E-16 puc = 7.986698224301345E-24 ud = 0
+ up = 0 lp = 1 eu = 1.67
+ vsat = 1.681183981233322E5 lvsat = -0.025321358592233 wvsat = -0.933385589369068
+ pvsat = 2.688877456410007E-7 a0 = 3.791647055136825 la0 = -7.975023877669317E-7
+ wa0 = -1.741884748655374E-5 pa0 = 4.584915005201252E-12 ags = 8.717042371324348
+ lags = -1.519692463411931E-6 wags = -2.331756237373842E-5 pags = 4.745590294303244E-12
+ b0 = 0 b1 = 0 keta = 0.384537234700585
+ lketa = -1.203363144642318E-7 wketa = -3.280860005181705E-6 pketa = 8.361199123424494E-13
+ a1 = 0 a2 = -0.102005265096319 la2 = 2.467164801091452E-7
+ wa2 = 7.827818857855366E-6 pa2 = -2.1410650140006E-12 rdsw = 531.92
+ rdswmin = 0 rdw = 0 rdwmin = 0
+ rsw = 0 rswmin = 0 prwb = -0.32348
+ prwg = 0.02 wr = 1 voff = -0.01976965408013
+ lvoff = -5.131355070755691E-8 wvoff = -8.265223302519349E-7 pvoff = 1.9058052789308E-13
+ voffl = 0 minv = 0 nfactor = 9.803997855166749
+ lnfactor = -1.916706519509882E-6 wnfactor = -5.250710559865244E-5 pnfactor = 1.268779195857879E-11
+ eta0 = 0.49 etab = -6.25E-4 dsub = 3.805262130725588
+ ldsub = -8.799610286543574E-7 wdsub = -1.938799659522906E-5 pdsub = 5.485227875859782E-12
+ cit = 1E-5 cdsc = 0 cdscb = 0
+ cdscd = 0 pclm = 1.233741351565131 lpclm = -8.241479669169022E-8
+ wpclm = -3.186471212346384E-6 ppclm = 4.700696622949763E-13 pdiblc1 = 0.926643593989753
+ lpdiblc1 = -1.144658025071164E-7 wpdiblc1 = -4.51759482872955E-6 ppdiblc1 = 9.81038929053836E-13
+ pdiblc2 = 5.066555977613928E-3 lpdiblc2 = 8.903203988209419E-10 wpdiblc2 = 1.024899240095717E-8
+ ppdiblc2 = -2.518619725367587E-15 pdiblcb = 0.924127787286042 lpdiblcb = -2.596054323784783E-7
+ wpdiblcb = -3.573565269432136E-6 ppdiblcb = 9.774415724950778E-13 drout = 0.448382312697603
+ ldrout = 1.114567315909902E-7 wdrout = 3.28759297554081E-7 pdrout = -6.507878801020743E-13
+ pscbe1 = 8E8 pscbe2 = -6.562293270276453E-8 lpscbe2 = 1.822270455286016E-14
+ wpscbe2 = 2.97004450724684E-13 ppscbe2 = -8.123665736221557E-20 pvag = 0
+ delta = 0.01 fprout = 0 pdits = 0
+ pditsl = 0 pditsd = 0 lambda = 0
+ vtl = 0 lc = 5E-9 xn = 3
+ alpha0 = 6.771515431421582E-8 lalpha0 = -3.522641393104549E-15 walpha0 = -3.368094749610824E-13
+ palpha0 = 1.754723493751268E-20 alpha1 = -2.490636E-10 walpha1 = 1.7387807368992E-15
+ beta0 = 43.083617851930036 lbeta0 = -1.895786144132959E-6 wbeta0 = -1.751256455500579E-4
+ pbeta0 = 1.065797079901992E-11 aigbacc = 0.43 bigbacc = 0.054
+ cigbacc = 0.075 nigbacc = 1 aigbinv = 0.35
+ bigbinv = 0.03 cigbinv = 6E-3 eigbinv = 1.1
+ nigbinv = 3 aigc = 0.43 bigc = 0.054
+ cigc = 0.075 aigsd = 0.43 bigsd = 0.054
+ cigsd = 0.075 dlcig = 0 nigc = 1
+ poxedge = 1 pigcd = 1 ntox = 1
+ toxref = 4.23E-9 agidl = 1E-10 bgidl = -1.259459367019385E9
+ lbgidl = 714.2032922469252 wbgidl = 1.432002699043101E4 pbgidl = -4.125721068821714E-3
+ cgidl = 2.846936635047339E3 lcgidl = -6.966381084181481E-4 wcgidl = -0.012686984145936
+ pcgidl = 3.470143903596286E-9 egidl = 0.1 noia = 1.2E41
+ noib = 2E25 noic = 0 em = 4.1E7
+ af = 1 ef = 0.88 kf = 0
+ lintnoi = -6E-8 tnoia = 1.5 tnoib = 3.5
+ ntnoi = 1 rnoia = 0.577 rnoib = 0.37
+ xpart = 0 cgso = {5.932020000000001E-11/sw_func_tox_lv_ratio} cgdo = {5.932020000000001E-11/sw_func_tox_lv_ratio}
+ cgbo = {0/sw_func_tox_lv_ratio} ckappas = 0.6 cf = 1.2E-11
+ clc = 1E-7 cle = 0.6 dlc = -2.56E-9
+ dwc = 0 vfbcv = -0.1446893 noff = 4
+ voffcv = -0.1375 acde = 0.552 moin = 14.504
+ cgsl = {7.513892E-12/sw_func_tox_lv_ratio} cgdl = {7.513892E-12/sw_func_tox_lv_ratio} ijthsrev = 0.1
+ ijthsfwd = 0.1 xjbvs = 1 bvs = 12.8
+ jss = 2.17E-5 jsws = 8.200000000000001E-10 cjs = {7.433E-04*sw_func_psd_nw_cj}
+ mjs = 0.34629 mjsws = 0.26859 cjsws = {9.2435E-11*sw_func_psd_nw_cj}
+ cjswgs = {2.4701E-10*sw_func_psd_nw_cj} mjswgs = 0.70393 pbs = 0.6587
+ pbsws = 0.7418 pbswgs = 1.3925 xrcrg1 = 12
+ xrcrg2 = 1 rbpb = 50 rbpd = 50
+ rbps = 50 rbdb = 50 rbsb = 50
+ gbmin = 1E-12 tnom = 30 ute = -1.648664104597762
+ lute = 4.215981144390197E-7 wute = 1.353430441014533E-5 pute = -3.592516941616917E-12
+ kt1 = -0.408712102875554 lkt1 = -3.738600878436729E-8 wkt1 = -1.93320832146553E-7
+ pkt1 = 1.455076524305839E-13 kt1l = 0 kt2 = 0.022027879404289
+ lkt2 = -1.528717673636084E-8 wkt2 = -1.229996659301633E-7 pkt2 = 2.503289201010684E-14
+ ua1 = 3.339621791377774E-9 lua1 = -6.028286397812046E-16 wua1 = 1.838248726260426E-15
+ pua1 = -3.741203807685219E-22 ub1 = -1.683862501667164E-18 lub1 = 3.570332028993013E-25
+ wub1 = -9.939761842480652E-24 pub1 = 2.022940330181662E-30 uc1 = -4.730024478824893E-10
+ luc1 = 9.436118260904423E-17 wuc1 = 1.469630745048587E-15 puc1 = -2.990992492322884E-22
+ at = 1.223245528711118E5 lat = -0.015639163246729 wat = -0.28899386780724
+ pat = 4.112219919744327E-8 prt = 0 njs = 1.2556
+ xtis = 2 tpb = 1.9551E-3 tpbsw = 1.4242E-4
+ tpbswg = 0 tcj = 1.2407E-3 tcjsw = 0
+ tcjswg = 2E-12 tvoff = 0 tvfbsdoff = 0
+ saref = 1.25E-6 sbref = 1.24E-6 wlod = 0
+ ku0 = 4.5E-8 kvsat = 0.4 kvth0 = 2.65E-8
+ tku0 = 0 llodku0 = 0 wlodku0 = 1
+ llodvth = 0 wlodvth = 1 lku0 = 0
+ wku0 = 2.5E-7 pku0 = 0 lkvth0 = 0
+ wkvth0 = 2.5E-7 pkvth0 = 0 stk2 = 0
+ lodk2 = 1 steta0 = 0 lodeta0 = 1

.model phighvt_model.16 pmos
+ level = 54 lmin = 1.5E-7 lmax = 1.8E-7 wmin = 5E-6
+ wmax = 7E-6 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 4.23E-9
+ toxm = 4.23E-9 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 9.999999999999999E22 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {9.364E-9+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {-1.176E-8-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = -5.722E-9 dwb = -1.7864E-8 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = -0.877491569526296 lvth0 = -3.951925469579792E-8
+ wvth0 = -5.674648089894993E-7 pvth0 = 9.84664936558579E-14 k1 = 3.262281482142357
+ lk1 = -4.182938401941419E-7 wk1 = -1.05559519015479E-5 pk1 = 1.831668773956592E-12
+ k2 = -0.957445547936116 lk2 = 1.455186604468349E-7 wk2 = 2.703361633289604E-6
+ pk2 = -4.479673842657395E-13 k3 = -13.778 k3b = 2
+ w0 = 0 lpe0 = 0 lpeb = 0
+ vbm = -3 dvtp0 = 0 dvtp1 = 0
+ dvt0 = 4.05 dvt1 = 0.3 dvt2 = 0.03
+ dvt0w = -4.254 dvt1w = 1.1472E6 dvt2w = -8.96E-3
+ vfbsdoff = 0 u0 = -0.027785008730557 lu0 = 5.17941908212632E-9
+ wu0 = 2.707227190470108E-7 pu0 = -4.697580620903732E-14 ua = -1.233806035044514E-8
+ lua = 1.687192865436441E-15 wua = 8.45196106389859E-14 pua = -1.46960141614235E-20
+ ub = 9.407210160382966E-18 lub = -1.252658273711252E-24 wub = -6.309052563155184E-23
+ pub = 1.10379819776269E-29 uc = 9.17809756524364E-11 luc = -1.431937962089076E-17
+ wuc = -1.532701133910101E-15 puc = 2.659543007560806E-22 ud = 0
+ up = 0 lp = 1 eu = 1.67
+ vsat = -1.070860696670717E5 lvsat = 0.03068825469247 wvsat = 2.329123782953512
+ pvsat = -3.950981618140908E-7 a0 = -7.606845263516146 la0 = 1.522318768925322E-6
+ wa0 = 3.466103882459442E-5 pa0 = -6.014383456843622E-12 ags = 1.25
+ b0 = 0 b1 = 0 keta = -0.048927596695228
+ lketa = -3.211755197855582E-8 wketa = 8.988813027210738E-9 pketa = 1.665698808605707E-13
+ a1 = 0 a2 = 4.914642377091403 la2 = -7.742716480289001E-7
+ wa2 = -1.826491066832914E-5 pa2 = 3.169327299168472E-12 rdsw = 531.92
+ rdswmin = 0 rdw = 0 rdwmin = 0
+ rsw = 0 rswmin = 0 prwb = -0.32348
+ prwg = 0.02 wr = 1 voff = -0.333684285051499
+ lvoff = 1.257435498773612E-8 wvoff = 7.455567746735372E-7 pvoff = -1.293690115413521E-13
+ voffl = 0 minv = 0 nfactor = -8.499985221144808
+ lnfactor = 1.808520116181047E-6 wnfactor = 6.671819423803473E-5 pnfactor = -1.157694106418379E-11
+ eta0 = 0.49 etab = -4.203850710414233E-3 letab = 7.283676752710774E-10
+ petab = -6.140467725170866E-22 dsub = -7.346928824596182 ldsub = 1.389732874572729E-6
+ wdsub = 5.131276029329208E-5 pdsub = -8.903790166092038E-12 cit = 1E-5
+ cdsc = 0 cdscb = 0 cdscd = 0
+ pclm = 0.841143932414844 lpclm = -2.513369946223719E-9 wpclm = -5.948031961391986E-6
+ ppclm = 1.032102505940737E-12 pdiblc1 = 1.384772990189269 lpdiblc1 = -2.07704297221642E-7
+ wpdiblc1 = 2.053934317026603E-6 ppdiblc1 = -3.56398682690456E-13 pdiblc2 = -0.145041614946102
+ lpdiblc2 = 3.144033534521563E-8 wpdiblc2 = -1.442482639749273E-8 ppdiblc2 = 2.502995876492938E-15
+ pdiblcb = -1.082831503667429 lpdiblcb = 1.488509225163722E-7 wpdiblcb = 8.338318962008299E-6
+ ppdiblcb = -1.446865106287679E-12 drout = 0.984014724506879 ldrout = 2.444823139566426E-9
+ wdrout = -1.946262626212889E-5 pdrout = 3.377154909004604E-12 pscbe1 = 7.9964807E8
+ pscbe2 = 1.083451920165837E-7 lpscbe2 = -1.71832881900216E-14 wpscbe2 = -6.930103850242611E-13
+ ppscbe2 = 1.202511620094098E-19 pvag = 0 delta = 0.01
+ fprout = 0 pdits = 0 pditsl = 0
+ pditsd = 0 lambda = 0 vtl = 0
+ lc = 5E-9 xn = 3 alpha0 = 3.413798270974879E-7
+ lalpha0 = -5.921887559795609E-14 walpha0 = -1.700007646885558E-12 palpha0 = 2.949853268875819E-19
+ alpha1 = -2.268047462399996E-9 lalpha1 = 4.109035956756473E-16 walpha1 = 1.179588851912416E-14
+ palpha1 = -2.046822575838423E-21 beta0 = 176.5375113683945 lbeta0 = -2.905632255260381E-5
+ wbeta0 = -8.327866861109275E-4 pbeta0 = 1.445051457739681E-10 aigbacc = 0.43
+ bigbacc = 0.054 cigbacc = 0.075 nigbacc = 1
+ aigbinv = 0.35 bigbinv = 0.03 cigbinv = 6E-3
+ eigbinv = 1.1 nigbinv = 3 aigc = 0.43
+ bigc = 0.054 cigc = 0.075 aigsd = 0.43
+ bigsd = 0.054 cigsd = 0.075 dlcig = 0
+ nigc = 1 poxedge = 1 pigcd = 1
+ ntox = 1 toxref = 4.23E-9 agidl = 1.563219430719998E-9
+ lagidl = -2.977944185401339E-16 wagidl = -8.045686225779966E-15 pagidl = 1.637458060670739E-21
+ bgidl = 9.478604062371315E9 lbgidl = -1.47120737690267E3 wbgidl = -4.037697252430641E4
+ pbgidl = 7.006212272417646E-3 cgidl = -5.642852148443778E3 lcgidl = 1.031203704797964E-3
+ wcgidl = 0.029602963007183 pcgidl = -5.136706141006364E-9 egidl = 0.1
+ noia = 1.2E41 noib = 2E25 noic = 0
+ em = 4.1E7 af = 1 ef = 0.88
+ kf = 0 lintnoi = -6E-8 tnoia = 1.5
+ tnoib = 3.5 ntnoi = 1 rnoia = 0.577
+ rnoib = 0.37 xpart = 0 cgso = {5.932020000000001E-11/sw_func_tox_lv_ratio}
+ cgdo = {5.932020000000001E-11/sw_func_tox_lv_ratio} cgbo = {0/sw_func_tox_lv_ratio} ckappas = 0.6
+ cf = 1.2E-11 clc = 1E-7 cle = 0.6
+ dlc = -2.56E-9 dwc = 0 vfbcv = -0.1446893
+ noff = 4 voffcv = -0.1375 acde = 0.552
+ moin = 14.504 cgsl = {7.513892E-12/sw_func_tox_lv_ratio} cgdl = {7.513892E-12/sw_func_tox_lv_ratio}
+ ijthsrev = 0.1 ijthsfwd = 0.1 xjbvs = 1
+ bvs = 12.8 jss = 2.17E-5 jsws = 8.200000000000001E-10
+ cjs = {7.433E-04*sw_func_psd_nw_cj} mjs = 0.34629 mjsws = 0.26859
+ cjsws = {9.2435E-11*sw_func_psd_nw_cj} cjswgs = {2.4701E-10*sw_func_psd_nw_cj} mjswgs = 0.70393
+ pbs = 0.6587 pbsws = 0.7418 pbswgs = 1.3925
+ xrcrg1 = 12 xrcrg2 = 1 rbpb = 50
+ rbpd = 50 rbps = 50 rbdb = 50
+ rbsb = 50 gbmin = 1E-12 tnom = 30
+ ute = 1.990551252029438 lute = -3.190549949417478E-7 wute = -2.089386815458044E-5
+ pute = 3.414304738756073E-12 kt1 = -0.25390834624 lkt1 = -6.889166933483522E-8
+ wkt1 = 1.52734499929225E-6 pkt1 = -2.046822575838413E-13 kt1l = 0
+ kt2 = -0.115281352 lkt2 = 1.265799803903998E-8 ua1 = 8.65085519999999E-10
+ lua1 = -9.921101783039981E-17 ub1 = 1.621275359999998E-19 lub1 = -1.866268956671996E-26
+ uc1 = 2.739337871999995E-10 luc1 = -5.76552799549439E-17 at = 1.342455673599998E5
+ lat = -0.018065328115507 wat = -1.595505204178703 pat = 3.070233863757634E-7
+ prt = 0 njs = 1.2556 xtis = 2
+ tpb = 1.9551E-3 tpbsw = 1.4242E-4 tpbswg = 0
+ tcj = 1.2407E-3 tcjsw = 0 tcjswg = 2E-12
+ tvoff = 0 tvfbsdoff = 0 saref = 1.1E-6
+ sbref = 1.1E-6 wlod = 0 ku0 = 4.5E-8
+ kvsat = 0.4 kvth0 = 2.65E-8 tku0 = 0
+ llodku0 = 0 wlodku0 = 1 llodvth = 0
+ wlodvth = 1 lku0 = 0 wku0 = 2.5E-7
+ pku0 = 0 lkvth0 = 0 wkvth0 = 2.5E-7
+ pkvth0 = 0 stk2 = 0 lodk2 = 1
+ steta0 = 0 lodeta0 = 1

.model phighvt_model.17 pmos
+ level = 54 lmin = 8E-6 lmax = 2.02E-5 wmin = 3E-6
+ wmax = 5E-6 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 4.23E-9
+ toxm = 4.23E-9 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 9.999999999999999E22 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {9.364E-9+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {-1.176E-8-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = -5.722E-9 dwb = -1.7864E-8 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = -1.138847253064 wvth0 = 1.750431586606173E-7
+ k1 = 0.357110682846 wk1 = 3.838972540719401E-7 k2 = 0.065118881721812
+ wk2 = -1.55112021691878E-7 k3 = -13.778 k3b = 2
+ w0 = 0 lpe0 = 0 lpeb = 0
+ vbm = -3 dvtp0 = 0 dvtp1 = 0
+ dvt0 = 4.05 dvt1 = 0.3 dvt2 = 0.03
+ dvt0w = -4.254 dvt1w = 1.1472E6 dvt2w = -8.96E-3
+ vfbsdoff = 0 u0 = 0.010287413997722 wu0 = -5.837841559230664E-9
+ ua = -1.63514826109372E-9 wua = 4.031285154165718E-15 ub = 2.39693498314628E-18
+ wub = -6.555952367877838E-24 uc = -3.536616325228398E-11 wuc = -2.201258753886169E-16
+ ud = 0 up = 0 lp = 1
+ eu = 1.67 vsat = 1.603125E5 a0 = 1.774979363198
+ wa0 = -3.959930081000292E-7 ags = 0.69029193838084 wags = -7.485422110281244E-7
+ b0 = 0 b1 = 0 keta = -0.078198667697108
+ wketa = 1.400085607824926E-7 a1 = 0 a2 = 0.8
+ rdsw = 531.92 rdswmin = 0 rdw = 0
+ rdwmin = 0 rsw = 0 rswmin = 0
+ prwb = -0.32348 prwg = 0.02 wr = 1
+ voff = -0.31074547418944 wvoff = 3.764537245550602E-7 voffl = 0
+ minv = 0 nfactor = -1.6110777650092 wnfactor = 1.228101212156531E-5
+ eta0 = 0.08 etab = -0.07 dsub = 0.56
+ cit = 1E-5 cdsc = 0 cdscb = 0
+ cdscd = 0 pclm = 0.3473505552473 wpclm = -8.562344069213488E-7
+ pdiblc1 = 0.39 pdiblc2 = -1.338660609284003E-5 wpdiblc2 = 8.955030236272135E-10
+ pdiblcb = -5.3533410154612E-3 wpdiblcb = 1.139745775749884E-8 drout = 0.56
+ pscbe1 = 6.1213795578692E8 wpscbe1 = 531.0290704864176 pscbe2 = 9.9692040994608E-9
+ wpscbe2 = -1.814606652851699E-15 pvag = 0 delta = 0.01
+ fprout = 0 pdits = 0 pditsl = 0
+ pditsd = 0 lambda = 0 vtl = 0
+ lc = 5E-9 xn = 3 alpha0 = 1.0328613626782E-9
+ walpha0 = -2.781113460434363E-15 alpha1 = -1.483780042970062E-10 walpha1 = 7.404823896265442E-16
+ beta0 = 3.5349445285428 wbeta0 = -1.594815144497851E-6 aigbacc = 0.43
+ bigbacc = 0.054 cigbacc = 0.075 nigbacc = 1
+ aigbinv = 0.35 bigbinv = 0.03 cigbinv = 6E-3
+ eigbinv = 1.1 nigbinv = 3 aigc = 0.43
+ bigc = 0.054 cigc = 0.075 aigsd = 0.43
+ bigsd = 0.054 cigsd = 0.075 dlcig = 0
+ nigc = 1 poxedge = 1 pigcd = 1
+ ntox = 1 toxref = 4.23E-9 agidl = 3.153236065612001E-11
+ wagidl = 3.410559347697678E-16 bgidl = 2.1218056173148E9 wbgidl = -3.344407676343329E3
+ cgidl = 300 egidl = 0.1 noia = 1.2E41
+ noib = 2E25 noic = 0 em = 4.1E7
+ af = 1 ef = 0.88 kf = 0
+ lintnoi = -6E-8 tnoia = 1.5 tnoib = 3.5
+ ntnoi = 1 rnoia = 0.577 rnoib = 0.37
+ xpart = 0 cgso = {5.932020000000001E-11/sw_func_tox_lv_ratio} cgdo = {5.932020000000001E-11/sw_func_tox_lv_ratio}
+ cgbo = {0/sw_func_tox_lv_ratio} ckappas = 0.6 cf = 1.2E-11
+ clc = 1E-7 cle = 0.6 dlc = -2.56E-9
+ dwc = 0 vfbcv = -0.1446893 noff = 4
+ voffcv = -0.1375 acde = 0.552 moin = 14.504
+ cgsl = {7.513892E-12/sw_func_tox_lv_ratio} cgdl = {7.513892E-12/sw_func_tox_lv_ratio} ijthsrev = 0.1
+ ijthsfwd = 0.1 xjbvs = 1 bvs = 12.8
+ jss = 2.17E-5 jsws = 8.200000000000001E-10 cjs = {7.433E-04*sw_func_psd_nw_cj}
+ mjs = 0.34629 mjsws = 0.26859 cjsws = {9.2435E-11*sw_func_psd_nw_cj}
+ cjswgs = {2.4701E-10*sw_func_psd_nw_cj} mjswgs = 0.70393 pbs = 0.6587
+ pbsws = 0.7418 pbswgs = 1.3925 xrcrg1 = 12
+ xrcrg2 = 1 rbpb = 50 rbpd = 50
+ rbps = 50 rbdb = 50 rbsb = 50
+ gbmin = 1E-12 tnom = 30 ute = -0.38209298144
+ wute = 1.562275412835917E-7 kt1 = -0.3961383314 wkt1 = -1.770925313504591E-7
+ kt1l = 0 kt2 = -0.037961 ua1 = 1.78304215E-9
+ wua1 = 2.134763218585201E-15 ub1 = 2.1268111264E-19 wub1 = -5.644982223642479E-24
+ uc1 = -3.3632933508E-10 wuc1 = 2.272353348812622E-15 at = 0
+ prt = 0 njs = 1.2556 xtis = 2
+ tpb = 1.9551E-3 tpbsw = 1.4242E-4 tpbswg = 0
+ tcj = 1.2407E-3 tcjsw = 0 tcjswg = 2E-12
+ tvoff = 0 tvfbsdoff = 0 saref = 3E-6
+ sbref = 3E-6 wlod = 0 ku0 = 4.5E-8
+ kvsat = 0.4 kvth0 = 2.65E-8 tku0 = 0
+ llodku0 = 0 wlodku0 = 1 llodvth = 0
+ wlodvth = 1 lku0 = 0 wku0 = 2.5E-7
+ pku0 = 0 lkvth0 = 0 wkvth0 = 2.5E-7
+ pkvth0 = 0 stk2 = 0 lodk2 = 1
+ steta0 = 0 lodeta0 = 1

.model phighvt_model.18 pmos
+ level = 54 lmin = 4E-6 lmax = 8E-6 wmin = 3E-6
+ wmax = 5E-6 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 4.23E-9
+ toxm = 4.23E-9 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 9.999999999999999E22 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {9.364E-9+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {-1.176E-8-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = -5.722E-9 dwb = -1.7864E-8 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = -1.128892739183389 lvth0 = -7.98702412113578E-8
+ wvth0 = 1.056808307118734E-7 pvth0 = 5.565300255433063E-13 k1 = 0.259828024674581
+ lk1 = 7.805493534915439E-7 wk1 = 5.729334777492635E-7 pk1 = -1.516735921399478E-12
+ k2 = 0.113120439505425 lk2 = -3.851414589079735E-7 wk2 = -2.734251945040983E-7
+ pk2 = 9.492881083223066E-13 k3 = -13.778 k3b = 2
+ w0 = 0 lpe0 = 0 lpeb = 0
+ vbm = -3 dvtp0 = 0 dvtp1 = 0
+ dvt0 = 4.05 dvt1 = 0.3 dvt2 = 0.03
+ dvt0w = -4.254 dvt1w = 1.1472E6 dvt2w = -8.96E-3
+ vfbsdoff = 0 u0 = 3.35485555283542E-3 lu0 = 5.562352133371961E-8
+ wu0 = 2.16580405929117E-8 pu0 = -2.206137603653573E-13 ua = -3.362611846966831E-9
+ lua = 1.386033863052462E-14 wua = 1.115043876719219E-14 pua = -5.712067139719018E-20
+ ub = 3.394594119475856E-18 lub = -8.00473803352308E-24 wub = -1.082353035648762E-23
+ pub = 3.424099734317034E-29 uc = 4.49011674518372E-11 luc = -6.440265332511302E-16
+ wuc = -5.590472244030001E-16 puc = 2.719342222243884E-21 ud = 0
+ up = 0 lp = 1 eu = 1.67
+ vsat = 2.31231338823365E5 lvsat = -0.569018721676046 wvsat = -0.028155072198585
+ pvsat = 2.259027848867907E-7 a0 = 1.605889794703494 la0 = 1.356693534607039E-6
+ wa0 = 2.02634521864218E-7 pa0 = -4.803099959218737E-12 ags = 0.387303700788649
+ lags = 2.431032184085698E-6 wags = 1.823564575970564E-7 pags = -7.469084085687511E-12
+ b0 = 0 b1 = 0 keta = -0.065127333179184
+ lketa = -1.048781139312577E-7 wketa = 8.23958808676366E-8 pketa = 4.622564895504454E-13
+ a1 = 0 a2 = 0.8 rdsw = 531.92
+ rdswmin = 0 rdw = 0 rdwmin = 0
+ rsw = 0 rswmin = 0 prwb = -0.32348
+ prwg = 0.02 wr = 1 voff = -0.346607885029239
+ lvoff = 2.877427706213459E-7 wvoff = 4.635599003656115E-7 pvoff = -6.988981437394738E-13
+ voffl = 0 minv = 0 nfactor = -2.982470789911596
+ lnfactor = 1.100339936316487E-5 wnfactor = 1.696179420965019E-5 pnfactor = -3.755634869939083E-11
+ eta0 = 0.08 etab = -0.07 dsub = 0.56
+ cit = 1E-5 cdsc = 0 cdscb = 0
+ cdscd = 0 pclm = 0.060210094259454 lpclm = 2.303877231545201E-6
+ wpclm = -1.717503472155395E-6 ppclm = 6.910409570286675E-12 pdiblc1 = 0.39
+ pdiblc2 = -2.43116125429506E-4 lpdiblc2 = 1.843239392988126E-9 wpdiblc2 = 1.796271605033355E-9
+ ppdiblc2 = -7.227334728283804E-15 pdiblcb = -7.019781344051118E-3 lpdiblcb = 1.337071730524778E-8
+ wpdiblcb = 1.962648360570135E-8 ppdiblcb = -6.60257534735698E-14 drout = 0.56
+ pscbe1 = 6.135808013854105E8 lpscbe1 = -11.576700516400082 wpscbe1 = 497.51802547759655
+ ppscbe1 = 2.688765398491752E-4 pscbe2 = 1.166373231927153E-8 lpscbe2 = -1.359608106221577E-14
+ wpscbe2 = -7.490527250730863E-15 ppscbe2 = 4.554086243549544E-20 pvag = 0
+ delta = 0.01 fprout = 0 pdits = 0
+ pditsl = 0 pditsd = 0 lambda = 0
+ vtl = 0 lc = 5E-9 xn = 3
+ alpha0 = 1.971207950168948E-9 lalpha0 = -7.528842611663765E-15 walpha0 = -5.57857986801608E-15
+ palpha0 = 2.244552767056006E-20 alpha1 = -3.982164712592787E-10 lalpha1 = 2.004583936441133E-15
+ walpha1 = 1.485318815704092E-15 palpha1 = -5.97620996136173E-21 beta0 = 2.172240540107943
+ lbeta0 = 1.093368270528684E-5 wbeta0 = -8.604491362038811E-6 pbeta0 = 5.624227732496426E-11
+ aigbacc = 0.43 bigbacc = 0.054 cigbacc = 0.075
+ nigbacc = 1 aigbinv = 0.35 bigbinv = 0.03
+ cigbinv = 6E-3 eigbinv = 1.1 nigbinv = 3
+ aigc = 0.43 bigc = 0.054 cigc = 0.075
+ aigsd = 0.43 bigsd = 0.054 cigsd = 0.075
+ dlcig = 0 nigc = 1 poxedge = 1
+ pigcd = 1 ntox = 1 toxref = 4.23E-9
+ agidl = -9.417951230436661E-9 lagidl = 7.581812058280474E-14 wagidl = 2.865027723748057E-14
+ pagidl = -2.271396033067262E-19 bgidl = 9.745385433076798E8 lbgidl = 9.205120313637612E3
+ wbgidl = -518.7374917101606 pbgidl = -0.022671821239808 cgidl = 300
+ egidl = -0.425564299150895 legidl = 4.216875665523186E-6 wegidl = 1.566850129258186E-6
+ pegidl = -1.257165334910564E-11 noia = 1.2E41 noib = 2E25
+ noic = 0 em = 4.1E7 af = 1
+ ef = 0.88 kf = 0 lintnoi = -6E-8
+ tnoia = 1.5 tnoib = 3.5 ntnoi = 1
+ rnoia = 0.577 rnoib = 0.37 xpart = 0
+ cgso = {5.932020000000001E-11/sw_func_tox_lv_ratio} cgdo = {5.932020000000001E-11/sw_func_tox_lv_ratio} cgbo = {0/sw_func_tox_lv_ratio}
+ ckappas = 0.6 cf = 1.2E-11 clc = 1E-7
+ cle = 0.6 dlc = -2.56E-9 dwc = 0
+ vfbcv = -0.1446893 noff = 4 voffcv = -0.1375
+ acde = 0.552 moin = 14.504 cgsl = {7.513892E-12/sw_func_tox_lv_ratio}
+ cgdl = {7.513892E-12/sw_func_tox_lv_ratio} ijthsrev = 0.1 ijthsfwd = 0.1
+ xjbvs = 1 bvs = 12.8 jss = 2.17E-5
+ jsws = 8.200000000000001E-10 cjs = {7.433E-04*sw_func_psd_nw_cj} mjs = 0.34629
+ mjsws = 0.26859 cjsws = {9.2435E-11*sw_func_psd_nw_cj} cjswgs = {2.4701E-10*sw_func_psd_nw_cj}
+ mjswgs = 0.70393 pbs = 0.6587 pbsws = 0.7418
+ pbswgs = 1.3925 xrcrg1 = 12 xrcrg2 = 1
+ rbpb = 50 rbpd = 50 rbps = 50
+ rbdb = 50 rbsb = 50 gbmin = 1E-12
+ tnom = 30 ute = 0.986634925619686 lute = -1.098201573685154E-5
+ wute = -2.446543065522239E-6 pute = 2.088338201911872E-11 kt1 = -0.304150270240784
+ lkt1 = -7.380680484721933E-7 wkt1 = -6.155183653136775E-7 pkt1 = 3.517718447320563E-12
+ kt1l = 0 kt2 = -0.0313322508 lkt2 = -5.318590178118399E-8
+ ua1 = 3.916344793042E-9 lua1 = -1.711659642250035E-14 wua1 = 4.282078844895683E-15
+ pua1 = -1.722902987401468E-20 ub1 = -1.318203049927283E-19 lub1 = 2.764114014404546E-24
+ wub1 = -1.2267303615184E-23 pub1 = 5.313432813146125E-29 uc1 = -7.356328498502703E-10
+ luc1 = 3.20381973682956E-15 wuc1 = 4.558068135316262E-15 puc1 = -1.833947830380769E-20
+ at = -1.896342590392288E5 lat = 1.521534270086433 wat = 0.027336261538422
+ pat = -2.193330411787607E-7 prt = 0 njs = 1.2556
+ xtis = 2 tpb = 1.9551E-3 tpbsw = 1.4242E-4
+ tpbswg = 0 tcj = 1.2407E-3 tcjsw = 0
+ tcjswg = 2E-12 tvoff = 0 tvfbsdoff = 0
+ saref = 3E-6 sbref = 3E-6 wlod = 0
+ ku0 = 4.5E-8 kvsat = 0.4 kvth0 = 2.65E-8
+ tku0 = 0 llodku0 = 0 wlodku0 = 1
+ llodvth = 0 wlodvth = 1 lku0 = 0
+ wku0 = 2.5E-7 pku0 = 0 lkvth0 = 0
+ wkvth0 = 2.5E-7 pkvth0 = 0 stk2 = 0
+ lodk2 = 1 steta0 = 0 lodeta0 = 1

.model phighvt_model.19 pmos
+ level = 54 lmin = 2E-6 lmax = 4E-6 wmin = 3E-6
+ wmax = 5E-6 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 4.23E-9
+ toxm = 4.23E-9 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 9.999999999999999E22 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {9.364E-9+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {-1.176E-8-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = -5.722E-9 dwb = -1.7864E-8 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = -1.198752661191896 lvth0 = 2.012125521883091E-7
+ wvth0 = 4.631530023899994E-7 pvth0 = -8.817664066470674E-13 k1 = 0.233709528374752
+ lk1 = 8.85637645723831E-7 wk1 = 1.089382744229986E-6 pk1 = -3.594679874069994E-12
+ k2 = 0.081445110326859 lk2 = -2.57695138451429E-7 wk2 = -2.815494144567874E-7
+ pk2 = 9.8197606978635E-13 k3 = -13.778 k3b = 2
+ w0 = 0 lpe0 = 0 lpeb = 0
+ vbm = -3 dvtp0 = 0 dvtp1 = 0
+ dvt0 = 4.05 dvt1 = 0.3 dvt2 = 0.03
+ dvt0w = -4.254 dvt1w = 1.1472E6 dvt2w = -8.96E-3
+ vfbsdoff = 0 u0 = 0.026302007623732 lu0 = -3.670480396657335E-8
+ wu0 = -6.805248403747314E-8 pu0 = 1.403383296954887E-13 ua = 2.071881724558466E-9
+ lua = -8.005454944378844E-15 wua = -1.052846122042275E-14 pua = 3.010481628097827E-20
+ ub = 4.022273773887978E-19 lub = 4.035109400599043E-24 wub = 1.380378206070421E-24
+ pub = -1.486167283645318E-29 uc = -2.08890378308692E-10 luc = 3.771088269472742E-16
+ wuc = 4.236329706628107E-16 puc = -1.234491196207307E-21 ud = 0
+ up = 0 lp = 1 eu = 1.67
+ vsat = 1.714936061623097E5 lvsat = -0.328662759559636 wvsat = -0.077511522699453
+ pvsat = 4.244894506060425E-7 a0 = 1.550031109801376 la0 = 1.58144207048441E-6
+ wa0 = 1.494793015481629E-6 pa0 = -1.000212550145826E-11 ags = 0.310963526580237
+ lags = 2.738188401816727E-6 wags = 6.344302743792833E-7 pags = -9.288012128987136E-12
+ b0 = 0 b1 = 0 keta = -0.036104208260345
+ lketa = -2.216532375047028E-7 wketa = -1.598034030502726E-8 pketa = 8.580751829630819E-13
+ a1 = 0 a2 = 0.8 rdsw = 531.92
+ rdswmin = 0 rdw = 0 rdwmin = 0
+ rsw = 0 rswmin = 0 prwb = -0.32348
+ prwg = 0.02 wr = 1 voff = -0.345344913198831
+ lvoff = 2.826611782022634E-7 wvoff = 6.058615844554928E-7 pvoff = -1.271451815708793E-12
+ voffl = 0 minv = 0 nfactor = -1.651034108538017
+ lnfactor = 5.646337246924648E-6 wnfactor = 1.443116292751527E-5 pnfactor = -2.737430312309531E-11
+ eta0 = 0.08 etab = -0.07 dsub = 0.56
+ cit = 1E-5 cdsc = 0 cdscb = 0
+ cdscd = 0 pclm = 0.620930693176364 lpclm = 4.780668739103634E-8
+ wpclm = 9.478412961103118E-7 ppclm = -3.813658411725762E-12 pdiblc1 = 0.39
+ pdiblc2 = 2.15E-4 pdiblcb = -0.041254876810969 lpdiblcb = 1.511163086183E-7
+ wpdiblcb = 1.827002065763629E-7 ppdiblcb = -7.221561393204861E-13 drout = 0.56
+ pscbe1 = 4.205172038329615E8 lpscbe1 = 765.2185455078293 wpscbe1 = 1.131341434694499E3
+ ppscbe1 = -2.281324623603218E-3 pscbe2 = -2.585559726001745E-9 lpscbe2 = 4.373623046778215E-14
+ wpscbe2 = 5.792334198723793E-14 ppscbe2 = -2.176531487208568E-19 pvag = 0
+ delta = 0.01 fprout = 0 pdits = 0
+ pditsl = 0 pditsd = 0 lambda = 0
+ vtl = 0 lc = 5E-9 xn = 3
+ alpha0 = -2.793179989910511E-3 lalpha0 = 1.123841595535674E-8 walpha0 = 8.327229593007693E-9
+ palpha0 = -3.350477481205831E-14 alpha1 = 3.51992587936E-10 lalpha1 = -1.013897217412255E-15
+ walpha1 = -7.512584466211347E-16 palpha1 = 3.022703385149068E-21 beta0 = -64.73634889427798
+ lbeta0 = 2.801417304663273E-4 wbeta0 = 2.095317689317954E-4 pbeta0 = -8.214333286924837E-10
+ aigbacc = 0.43 bigbacc = 0.054 cigbacc = 0.075
+ nigbacc = 1 aigbinv = 0.35 bigbinv = 0.03
+ cigbinv = 6E-3 eigbinv = 1.1 nigbinv = 3
+ aigc = 0.43 bigc = 0.054 cigc = 0.075
+ aigsd = 0.43 bigsd = 0.054 cigsd = 0.075
+ dlcig = 0 nigc = 1 poxedge = 1
+ pigcd = 1 ntox = 1 toxref = 4.23E-9
+ agidl = 1.886122672405911E-8 lagidl = -3.796371750066811E-14 wagidl = -5.593231991808919E-14
+ pagidl = 1.131801680006518E-19 bgidl = 5.092119604706383E9 lbgidl = -7.362049438521299E3
+ wbgidl = -1.17762299311407E4 pbgidl = 0.02262292474009 cgidl = 300
+ egidl = 1.151128598301789 legidl = -2.126979741235637E-6 wegidl = -3.133700258516373E-6
+ pegidl = 6.341105147113051E-12 noia = 1.2E41 noib = 2E25
+ noic = 0 em = 4.1E7 af = 1
+ ef = 0.88 kf = 0 lintnoi = -6E-8
+ tnoia = 1.5 tnoib = 3.5 ntnoi = 1
+ rnoia = 0.577 rnoib = 0.37 xpart = 0
+ cgso = {5.932020000000001E-11/sw_func_tox_lv_ratio} cgdo = {5.932020000000001E-11/sw_func_tox_lv_ratio} cgbo = {0/sw_func_tox_lv_ratio}
+ ckappas = 0.6 cf = 1.2E-11 clc = 1E-7
+ cle = 0.6 dlc = -2.56E-9 dwc = 0
+ vfbcv = -0.1446893 noff = 4 voffcv = -0.1375
+ acde = 0.552 moin = 14.504 cgsl = {7.513892E-12/sw_func_tox_lv_ratio}
+ cgdl = {7.513892E-12/sw_func_tox_lv_ratio} ijthsrev = 0.1 ijthsfwd = 0.1
+ xjbvs = 1 bvs = 12.8 jss = 2.17E-5
+ jsws = 8.200000000000001E-10 cjs = {7.433E-04*sw_func_psd_nw_cj} mjs = 0.34629
+ mjsws = 0.26859 cjsws = {9.2435E-11*sw_func_psd_nw_cj} cjswgs = {2.4701E-10*sw_func_psd_nw_cj}
+ mjswgs = 0.70393 pbs = 0.6587 pbsws = 0.7418
+ pbswgs = 1.3925 xrcrg1 = 12 xrcrg2 = 1
+ rbpb = 50 rbpd = 50 rbps = 50
+ rbdb = 50 rbsb = 50 gbmin = 1E-12
+ tnom = 30 ute = -3.335977104739992 lute = 6.410100219541237E-6
+ wute = 5.01254599553038E-6 pute = -9.12841199980771E-12 kt1 = -0.557404991899112
+ lkt1 = 2.809073892145237E-7 wkt1 = 6.407332863058682E-7 pkt1 = -1.536835198003712E-12
+ kt1l = 0 kt2 = -0.039709935389811 lkt2 = -1.947812028038877E-8
+ wkt2 = -1.154954685497427E-9 pkt2 = 4.646983276192608E-15 ua1 = -2.370081736365121E-9
+ lua1 = 8.176966447099789E-15 wua1 = -2.84897336685104E-15 pua1 = 1.14629013209925E-20
+ ub1 = 2.114256972979399E-18 lub1 = -6.273022835061867E-24 wub1 = 3.267379226568917E-24
+ pub1 = -9.369778975988462E-30 uc1 = 2.798421020968221E-11 luc1 = 1.313912233371395E-16
+ wuc1 = 1.92976162863132E-16 puc1 = -7.764434508030689E-22 at = 3.718000332619278E5
+ lat = -0.737407833673117 wat = -0.28484354422028 pat = 1.036728650887492E-6
+ prt = 0 njs = 1.2556 xtis = 2
+ tpb = 1.9551E-3 tpbsw = 1.4242E-4 tpbswg = 0
+ tcj = 1.2407E-3 tcjsw = 0 tcjswg = 2E-12
+ tvoff = 0 tvfbsdoff = 0 saref = 3E-6
+ sbref = 3E-6 wlod = 0 ku0 = 4.5E-8
+ kvsat = 0.4 kvth0 = 2.65E-8 tku0 = 0
+ llodku0 = 0 wlodku0 = 1 llodvth = 0
+ wlodvth = 1 lku0 = 0 wku0 = 2.5E-7
+ pku0 = 0 lkvth0 = 0 wkvth0 = 2.5E-7
+ pkvth0 = 0 stk2 = 0 lodk2 = 1
+ steta0 = 0 lodeta0 = 1

.model phighvt_model.20 pmos
+ level = 54 lmin = 1E-6 lmax = 2E-6 wmin = 3E-6
+ wmax = 5E-6 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 4.23E-9
+ toxm = 4.23E-9 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 9.999999999999999E22 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {9.364E-9+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {-1.176E-8-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = -5.722E-9 dwb = -1.7864E-8 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = -1.09990029888414 lvth0 = 1.182820011319643E-9
+ wvth0 = -5.632892445466352E-9 pvth0 = 6.68312272703942E-14 k1 = 0.919597349802956
+ lk1 = -5.022700786925675E-7 wk1 = -1.453676531849636E-6 pk1 = 1.551251432262641E-12
+ k2 = -0.128537045035596 lk2 = 1.672079525676043E-7 wk2 = 4.615143665494059E-7
+ pk2 = -5.21628352355302E-13 k3 = -13.778 k3b = 2
+ w0 = 0 lpe0 = 0 lpeb = 0
+ vbm = -3 dvtp0 = 0 dvtp1 = 0
+ dvt0 = 4.05 dvt1 = 0.3 dvt2 = 0.03
+ dvt0w = -4.254 dvt1w = 1.1472E6 dvt2w = -8.96E-3
+ vfbsdoff = 0 u0 = 4.196184473355249E-3 lu0 = 8.026771294676583E-9
+ wu0 = 1.331808242005335E-8 pu0 = -2.43166389426453E-14 ua = -3.413120761001292E-9
+ lua = 3.093557285201038E-15 wua = 1.001561822621936E-14 pua = -1.146653936089096E-20
+ ub = 3.82843620793236E-18 lub = -2.897892692182465E-24 wub = -1.185315737213492E-23
+ pub = 1.191665107675688E-29 uc = 2.528989017531772E-11 luc = -9.675962993548915E-17
+ wuc = -4.412533190470003E-16 puc = 5.156235087462895E-22 ud = 0
+ up = 0 lp = 1 eu = 1.67
+ vsat = -6.532160437775103E4 lvsat = 0.150537555272387 wvsat = 0.313767161057706
+ pvsat = -3.672707915502444E-7 a0 = 3.653392562778307 la0 = -2.674751896843469E-6
+ wa0 = -7.462914825530105E-6 pa0 = 8.123975468985798E-12 ags = 2.729288283248497
+ lags = -2.15534010979663E-6 wags = -7.869667600247347E-6 pags = 7.920200002277339E-12
+ b0 = 0 b1 = 0 keta = -0.282874532065846
+ lketa = 2.776914481222053E-7 wketa = 8.361277156542628E-7 pketa = -8.661825104316608E-13
+ a1 = 0 a2 = 0.8 rdsw = 531.92
+ rdswmin = 0 rdw = 0 rdwmin = 0
+ rsw = 0 rswmin = 0 prwb = -0.32348
+ prwg = 0.02 wr = 1 voff = -0.204922755026482
+ lvoff = -1.485867302649686E-9 wvoff = -5.052876758020274E-8 pvoff = 5.676718944247749E-14
+ voffl = 0 minv = 0 nfactor = 0.84430787928009
+ lnfactor = 5.969628277349521E-7 wnfactor = 7.370578731449484E-7 pnfactor = 3.35992336524113E-13
+ eta0 = -0.064825330875719 leta0 = 2.93056953533635E-7 weta0 = 7.633953140354877E-9
+ peta0 = -1.54474568585709E-14 etab = -0.638113720015354 letab = 1.14958947472547E-6
+ wetab = 4.021247287905655E-6 petab = -8.13707431202285E-12 dsub = 0.071869155067831
+ ldsub = 9.877425273371427E-7 wdsub = 9.358161955303733E-7 pdsub = -1.893642787979621E-12
+ cit = 1E-5 cdsc = 0 cdscb = 0
+ cdscd = 0 pclm = 0.714455289636076 lpclm = -1.414422040371202E-7
+ wpclm = -2.037722091235141E-6 ppclm = 2.227688813835508E-12 pdiblc1 = 0.376959920135301
+ lpdiblc1 = 2.638686240781491E-8 wpdiblc1 = 9.690198789407784E-8 ppdiblc1 = -1.960831105434244E-13
+ pdiblc2 = -5.056799999999948E-6 lpdiblc2 = 4.452893359359999E-10 pdiblcb = 0.093224240293769
+ lpdiblcb = -1.21004874425478E-7 wpdiblcb = -3.524586173090842E-7 ppdiblcb = 3.607484439881938E-13
+ drout = 0.853068846472728 ldrout = -5.930306722144937E-7 wdrout = -2.186985988471022E-6
+ pdrout = 4.425409887390881E-12 pscbe1 = 8E8 pscbe2 = 2.919713529603096E-8
+ lpscbe2 = -2.057668856320148E-14 wpscbe2 = -1.010373882907258E-13 ppscbe2 = 1.040070682112084E-19
+ pvag = 0 delta = 0.01 fprout = 0
+ pdits = 0 pditsl = 0 pditsd = 0
+ lambda = 0 vtl = 0 lc = 5E-9
+ xn = 3 alpha0 = 5.550299318422883E-3 lalpha0 = -5.644781294642048E-9
+ walpha0 = -1.654695165150603E-8 palpha0 = 1.682862841984009E-14 alpha1 = -1.490636E-10
+ walpha1 = 7.425263368992002E-16 beta0 = 91.08816238495922 lbeta0 = -3.517228459743473E-5
+ wbeta0 = -2.514104107699628E-4 pbeta0 = 1.112923907776182E-10 aigbacc = 0.43
+ bigbacc = 0.054 cigbacc = 0.075 nigbacc = 1
+ aigbinv = 0.35 bigbinv = 0.03 cigbinv = 6E-3
+ eigbinv = 1.1 nigbinv = 3 aigc = 0.43
+ bigc = 0.054 cigc = 0.075 aigsd = 0.43
+ bigsd = 0.054 cigsd = 0.075 dlcig = 0
+ nigc = 1 poxedge = 1 pigcd = 1
+ ntox = 1 toxref = 4.23E-9 agidl = 1E-10
+ bgidl = 1.263660398696014E9 lbgidl = 384.9143340248017 wbgidl = 17.771176861437926
+ pbgidl = -1.24247238197484E-3 cgidl = 300 egidl = 0.1
+ noia = 1.2E41 noib = 2E25 noic = 0
+ em = 4.1E7 af = 1 ef = 0.88
+ kf = 0 lintnoi = -6E-8 tnoia = 1.5
+ tnoib = 3.5 ntnoi = 1 rnoia = 0.577
+ rnoib = 0.37 xpart = 0 cgso = {5.932020000000001E-11/sw_func_tox_lv_ratio}
+ cgdo = {5.932020000000001E-11/sw_func_tox_lv_ratio} cgbo = {0/sw_func_tox_lv_ratio} ckappas = 0.6
+ cf = 1.2E-11 clc = 1E-7 cle = 0.6
+ dlc = -2.56E-9 dwc = 0 vfbcv = -0.1446893
+ noff = 4 voffcv = -0.1375 acde = 0.552
+ moin = 14.504 cgsl = {7.513892E-12/sw_func_tox_lv_ratio} cgdl = {7.513892E-12/sw_func_tox_lv_ratio}
+ ijthsrev = 0.1 ijthsfwd = 0.1 xjbvs = 1
+ bvs = 12.8 jss = 2.17E-5 jsws = 8.200000000000001E-10
+ cjs = {7.433E-04*sw_func_psd_nw_cj} mjs = 0.34629 mjsws = 0.26859
+ cjsws = {9.2435E-11*sw_func_psd_nw_cj} cjswgs = {2.4701E-10*sw_func_psd_nw_cj} mjswgs = 0.70393
+ pbs = 0.6587 pbsws = 0.7418 pbswgs = 1.3925
+ xrcrg1 = 12 xrcrg2 = 1 rbpb = 50
+ rbpd = 50 rbps = 50 rbdb = 50
+ rbsb = 50 gbmin = 1E-12 tnom = 30
+ ute = 3.315259226562248 lute = -7.048809521575472E-6 wute = -9.88368950489169E-6
+ pute = 2.101441846000635E-11 kt1 = -0.34386735383896 lkt1 = -1.511902921529557E-7
+ wkt1 = -2.984378560583061E-7 pkt1 = 3.635963919930422E-13 kt1l = 0
+ kt2 = -0.038134316271672 lkt2 = -2.266641707832483E-8 wkt2 = -6.759402200144063E-8
+ pkt2 = 1.3908776477135E-13 ua1 = 8.040603263453486E-9 lua1 = -1.288926286373316E-14
+ wua1 = -1.552927349646055E-14 pua1 = 3.712174223925993E-20 ub1 = -4.88719248169956E-18
+ lub1 = 7.894550165470098E-24 wub1 = 1.000868159539859E-23 pub1 = -2.301093914536268E-29
+ uc1 = -4.461870144926965E-11 luc1 = 2.783046671372617E-16 wuc1 = 6.016478023359909E-16
+ puc1 = -1.603398686709188E-21 at = -1.063506057923998E5 lat = 0.230139547466096
+ wat = 0.50867744167029 pat = -5.689769344817948E-7 prt = 0
+ njs = 1.2556 xtis = 2 tpb = 1.9551E-3
+ tpbsw = 1.4242E-4 tpbswg = 0 tcj = 1.2407E-3
+ tcjsw = 0 tcjswg = 2E-12 tvoff = 0
+ tvfbsdoff = 0 saref = 3E-6 sbref = 3E-6
+ wlod = 0 ku0 = 4.5E-8 kvsat = 0.4
+ kvth0 = 2.65E-8 tku0 = 0 llodku0 = 0
+ wlodku0 = 1 llodvth = 0 wlodvth = 1
+ lku0 = 0 wku0 = 2.5E-7 pku0 = 0
+ lkvth0 = 0 wkvth0 = 2.5E-7 pkvth0 = 0
+ stk2 = 0 lodk2 = 1 steta0 = 0
+ lodeta0 = 1

.model phighvt_model.21 pmos
+ level = 54 lmin = 5E-7 lmax = 1E-6 wmin = 3E-6
+ wmax = 5E-6 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 4.23E-9
+ toxm = 4.23E-9 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 9.999999999999999E22 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {9.364E-9+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {-1.176E-8-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = -5.722E-9 dwb = -1.7864E-8 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = -1.127108471321232 lvth0 = 2.903092866413126E-8
+ wvth0 = 4.968224274318806E-8 pvth0 = 1.021508010210265E-14 k1 = 0.505595937533109
+ lk1 = -7.853135320613426E-8 wk1 = -5.396698085289807E-7 pk1 = 6.157472708094848E-13
+ k2 = 0.010395302538254 lk2 = 2.500791617881749E-8 wk2 = 1.288418682694905E-7
+ pk2 = -1.811313969158431E-13 k3 = -13.778 k3b = 2
+ w0 = 0 lpe0 = 0 lpeb = 0
+ vbm = -3 dvtp0 = 0 dvtp1 = 0
+ dvt0 = 4.05 dvt1 = 0.3 dvt2 = 0.03
+ dvt0w = -4.254 dvt1w = 1.1472E6 dvt2w = -8.96E-3
+ vfbsdoff = 0 u0 = 0.016106122782316 lu0 = -4.163288763311263E-9
+ wu0 = -1.399418618276467E-8 pu0 = 3.638014217711E-15 ua = 6.84894407709946E-10
+ lua = -1.100843200278288E-15 wua = -2.840566974135982E-15 pua = 1.692023315376736E-21
+ ub = 2.107514271840762E-19 lub = 8.048800346090174E-25 wub = 1.71503846394938E-24
+ pub = -1.970668725392115E-30 uc = -1.636235744255624E-10 luc = 9.65970793528036E-17
+ wuc = 2.929718161143595E-16 puc = -2.358706015940654E-22 ud = 0
+ up = 0 lp = 1 eu = 1.67
+ vsat = -5.659486771128548E4 lvsat = 0.141605565759527 wvsat = 0.404910496543298
+ pvsat = -4.605578182864577E-7 a0 = 0.662577074281071 la0 = 3.864075719432216E-7
+ wa0 = 1.658335795314105E-6 pa0 = -1.211806966460666E-12 ags = 0.360830570398623
+ lags = 2.688237284594728E-7 wags = -1.450855619051794E-6 pags = 1.350417563284068E-12
+ b0 = 0 b1 = 0 keta = -0.012880420025824
+ lketa = 1.347074567001614E-9 wketa = 9.363987754214418E-8 pketa = -1.062313583671452E-13
+ a1 = 0 a2 = 1.030558658117889 la2 = -2.35981397756822E-7
+ wa2 = -1.311660278780436E-6 pa2 = 1.342510528537352E-12 rdsw = 531.92
+ rdswmin = 0 rdw = 0 rdwmin = 0
+ rsw = 0 rswmin = 0 prwb = -0.32348
+ prwg = 0.02 wr = 1 voff = -0.141653394425584
+ lvoff = -6.624332326488102E-8 wvoff = -2.354536005058196E-7 pvoff = 2.460414544385048E-13
+ voffl = 0 minv = 0 nfactor = 4.585070822823565
+ lnfactor = -3.231782860240664E-6 wnfactor = -1.206196041465491E-5 pnfactor = 1.343604353445302E-11
+ eta0 = 0.429844404156609 leta0 = -2.132474136666538E-7 weta0 = -1.840075693414035E-7
+ peta0 = 1.807014742319584E-13 etab = 0.992480562011706 letab = -5.193563848148669E-7
+ wetab = -8.03958074738172E-6 petab = 4.207424398654482E-12 dsub = 1.075564089864338
+ ldsub = -3.955931232577854E-8 wdsub = -1.871632391060747E-6 pdsub = 9.798369893681223E-13
+ cit = 1E-5 cdsc = 0 cdscb = 0
+ cdscd = 0 pclm = 0.641929124512144 lpclm = -6.721022350947316E-8
+ wpclm = -3.281358506940606E-7 ppclm = 4.778931049169013E-13 pdiblc1 = 1.351757862964943
+ lpdiblc1 = -9.713383280371797E-7 wpdiblc1 = -4.887435444745398E-6 ppdiblc1 = 4.905485938511731E-12
+ pdiblc2 = -1.719686926880322E-3 lpdiblc2 = 2.200247563400546E-9 wpdiblc2 = 4.574733599695639E-9
+ ppdiblc2 = -4.68233133396048E-15 pdiblcb = 0.01349796040417 lpdiblcb = -3.940343243287577E-8
+ wpdiblcb = -1.917688122183992E-7 ppdiblcb = 1.962792146817759E-13 drout = 0.234076961151461
+ ldrout = 4.051990224952861E-8 wdrout = 2.314556472264507E-6 pdrout = -1.820088520211457E-13
+ pscbe1 = 7.863501316862353E8 lpscbe1 = 13.970913216504407 wpscbe1 = 67.99370683504313
+ ppscbe1 = -6.959291881980333E-5 pscbe2 = 8.798412926354168E-9 lpscbe2 = 3.018117566101133E-16
+ wpscbe2 = 1.615384158814658E-15 ppscbe2 = -1.060097446345214E-21 pvag = 0
+ delta = 0.01 fprout = 0 pdits = 0
+ pditsl = 0 pditsd = 0 lambda = 0
+ vtl = 0 lc = 5E-9 xn = 3
+ alpha0 = 7.212202279628058E-5 lalpha0 = -3.775726902230881E-11 walpha0 = -2.15015069018713E-10
+ palpha0 = 1.125646889326766E-16 alpha1 = -4.098431517440001E-10 lalpha1 = 2.669130868010189E-16
+ walpha1 = 1.519981112686139E-15 palpha1 = -7.957405121134473E-22 beta0 = 106.74164890204952
+ lbeta0 = -5.119394111740698E-5 wbeta0 = -2.930866800420434E-4 pbeta0 = 1.53948885902978E-10
+ aigbacc = 0.43 bigbacc = 0.054 cigbacc = 0.075
+ nigbacc = 1 aigbinv = 0.35 bigbinv = 0.03
+ cigbinv = 6E-3 eigbinv = 1.1 nigbinv = 3
+ aigc = 0.43 bigc = 0.054 cigc = 0.075
+ aigsd = 0.43 bigsd = 0.054 cigsd = 0.075
+ dlcig = 0 nigc = 1 poxedge = 1
+ pigcd = 1 ntox = 1 toxref = 4.23E-9
+ agidl = 1E-10 bgidl = 2.185674947296288E9 lbgidl = -558.7859967585503
+ wbgidl = -2.689980933589826E3 pbgidl = 1.528966058114238E-3 cgidl = 300
+ egidl = 0.1 noia = 1.2E41 noib = 2E25
+ noic = 0 em = 4.1E7 af = 1
+ ef = 0.88 kf = 0 lintnoi = -6E-8
+ tnoia = 1.5 tnoib = 3.5 ntnoi = 1
+ rnoia = 0.577 rnoib = 0.37 xpart = 0
+ cgso = {5.932020000000001E-11/sw_func_tox_lv_ratio} cgdo = {5.932020000000001E-11/sw_func_tox_lv_ratio} cgbo = {0/sw_func_tox_lv_ratio}
+ ckappas = 0.6 cf = 1.2E-11 clc = 1E-7
+ cle = 0.6 dlc = -2.56E-9 dwc = 0
+ vfbcv = -0.1446893 noff = 4 voffcv = -0.1375
+ acde = 0.552 moin = 14.504 cgsl = {7.513892E-12/sw_func_tox_lv_ratio}
+ cgdl = {7.513892E-12/sw_func_tox_lv_ratio} ijthsrev = 0.1 ijthsfwd = 0.1
+ xjbvs = 1 bvs = 12.8 jss = 2.17E-5
+ jsws = 8.200000000000001E-10 cjs = {7.433E-04*sw_func_psd_nw_cj} mjs = 0.34629
+ mjsws = 0.26859 cjsws = {9.2435E-11*sw_func_psd_nw_cj} cjswgs = {2.4701E-10*sw_func_psd_nw_cj}
+ mjswgs = 0.70393 pbs = 0.6587 pbsws = 0.7418
+ pbswgs = 1.3925 xrcrg1 = 12 xrcrg2 = 1
+ rbpb = 50 rbpd = 50 rbps = 50
+ rbdb = 50 rbsb = 50 gbmin = 1E-12
+ tnom = 30 ute = -7.05550839943936 lute = 3.565878558989694E-6
+ wute = 2.109681985771098E-5 pute = -1.069475248280473E-11 kt1 = -0.492010162014811
+ lkt1 = 4.36834871191674E-10 wkt1 = 1.170410050191037E-7 pkt1 = -6.165453189690834E-14
+ kt1l = 0 kt2 = -0.108428984297315 lkt2 = 4.928158153928106E-8
+ wkt2 = 2.437762368488466E-7 pkt2 = -1.79605922567096E-13 ua1 = -1.250648106804874E-8
+ lua1 = 8.141088891245993E-15 wua1 = 4.524161583152145E-14 pua1 = -2.50784784057162E-20
+ ub1 = 8.19222621118286E-18 lub1 = -5.492496455068916E-24 wub1 = -2.748667311445742E-23
+ pub1 = 1.536630630726914E-29 uc1 = 8.301520090836697E-10 luc1 = -6.170406505074121E-16
+ wuc1 = -2.843773664579409E-15 puc1 = 1.923059093108062E-21 at = 1.651193587984999E5
+ lat = -0.047715390691981 wat = 0.02499309909606 pat = -7.391633617021811E-8
+ prt = 0 njs = 1.2556 xtis = 2
+ tpb = 1.9551E-3 tpbsw = 1.4242E-4 tpbswg = 0
+ tcj = 1.2407E-3 tcjsw = 0 tcjswg = 2E-12
+ tvoff = 0 tvfbsdoff = 0 saref = 2.75E-6
+ sbref = 2.74E-6 wlod = 0 ku0 = 4.5E-8
+ kvsat = 0.4 kvth0 = 2.65E-8 tku0 = 0
+ llodku0 = 0 wlodku0 = 1 llodvth = 0
+ wlodvth = 1 lku0 = 0 wku0 = 2.5E-7
+ pku0 = 0 lkvth0 = 0 wkvth0 = 2.5E-7
+ pkvth0 = 0 stk2 = 0 lodk2 = 1
+ steta0 = 0 lodeta0 = 1

.model phighvt_model.22 pmos
+ level = 54 lmin = 2.5E-7 lmax = 5E-7 wmin = 3E-6
+ wmax = 5E-6 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 4.23E-9
+ toxm = 4.23E-9 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 9.999999999999999E22 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {9.364E-9+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {-1.176E-8-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = -5.722E-9 dwb = -1.7864E-8 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = -1.085306390479894 lvth0 = 7.146703302074078E-9
+ wvth0 = 1.290736862702044E-7 pvth0 = -3.134792841316096E-14 k1 = -0.225901036682333
+ lk1 = 3.044219427351342E-7 wk1 = 2.023433283722631E-6 pk1 = -7.260884600460795E-13
+ k2 = 0.271492754775305 lk2 = -1.116818220163233E-7 wk2 = -7.479847938861925E-7
+ pk2 = 2.779048972559E-13 k3 = -13.778 k3b = 2
+ w0 = 0 lpe0 = 0 lpeb = 0
+ vbm = -3 dvtp0 = 0 dvtp1 = 0
+ dvt0 = 4.05 dvt1 = 0.3 dvt2 = 0.03
+ dvt0w = -4.254 dvt1w = 1.1472E6 dvt2w = -8.96E-3
+ vfbsdoff = 0 u0 = 0.012915521827708 lu0 = -2.492945351554599E-9
+ wu0 = -2.03915591854953E-8 pu0 = 6.987166932100539E-15 ua = -4.73494776124246E-10
+ lua = -4.944032947574117E-16 wua = -1.691183894243218E-15 pua = 1.090298285391277E-21
+ ub = 1.453488264025482E-18 lub = 1.54282445785805E-25 wub = -2.303209760675558E-24
+ pub = 1.329645851635324E-31 uc = 4.882544602412327E-11 luc = -1.462423183301579E-17
+ wuc = -2.814205802151236E-16 puc = 6.483530573234556E-23 ud = 0
+ up = 0 lp = 1 eu = 1.67
+ vsat = 3.470113358188638E5 lvsat = -0.069690353912577 wvsat = -0.957774491165159
+ pvsat = 2.528350264786738E-7 a0 = 2.170576840538738 la0 = -4.030604656879925E-7
+ wa0 = -1.631984284321709E-6 pa0 = 5.107414016302751E-13 ags = 0.171344852637824
+ lags = 3.680232914216062E-7 wags = -6.800044312901697E-8 pags = 6.264652215849759E-13
+ b0 = 0 b1 = 0 keta = 0.142226274979962
+ lketa = -7.985438240242725E-8 wketa = -4.977592542588856E-7 pketa = 2.033779151133299E-13
+ a1 = 0 a2 = 0.338882683764222 la2 = 1.261248083368101E-7
+ wa2 = 2.623320557560872E-6 pa2 = -7.175306389040495E-13 rdsw = 531.92
+ rdswmin = 0 rdw = 0 rdwmin = 0
+ rsw = 0 rswmin = 0 prwb = -0.32348
+ prwg = 0.02 wr = 1 voff = -0.303393656188358
+ lvoff = 1.843093857316651E-8 wvoff = 4.770063628347197E-7 pvoff = -1.269455855695343E-13
+ voffl = 0 minv = 0 nfactor = -4.719699832915854
+ lnfactor = 1.639450673452036E-6 wnfactor = 2.688516906291783E-5 pnfactor = -6.953557689645857E-12
+ eta0 = -0.488960284810342 leta0 = 2.677652171013248E-7 weta0 = 3.374793261213875E-7
+ peta0 = -9.230734528072189E-14 etab = 1.591956038006531E-3 letab = -6.063818155155463E-10
+ wetab = -5.827656859183461E-9 petab = 1.59398070412386E-15 dsub = 1.082878138297357
+ ldsub = -4.338836296143253E-8 wdsub = 1.103143859707141E-6 pdsub = -5.775178734338823E-13
+ cit = 1E-5 cdsc = 0 cdscb = 0
+ cdscd = 0 pclm = 0.379022936503842 lpclm = 7.042642403663304E-8
+ wpclm = 1.217641748257651E-6 ppclm = -3.313523836862989E-13 pdiblc1 = -1.314805471292176
+ lpdiblc1 = 4.246609087131069E-7 wpdiblc1 = 8.93216870439498E-6 ppdiblc1 = -2.329353225646239E-12
+ pdiblc2 = -4.97178375977579E-3 lpdiblc2 = 3.902785297357982E-9 wpdiblc2 = -4.972626522170731E-9
+ ppdiblc2 = 3.159026370390013E-16 pdiblcb = -0.101995920808339 lpdiblcb = 2.105992425949699E-8
+ wpdiblcb = 3.835376244367983E-7 ppdiblcb = -1.049052110359531E-13 drout = 0.156752779744921
+ ldrout = 8.100065769948097E-8 wdrout = 4.166098876794349E-6 pdrout = -1.151328331640609E-12
+ pscbe1 = 8.270594434998902E8 lpscbe1 = -7.341225704180136 wpscbe1 = -134.79044824158458
+ ppscbe1 = 3.656864204591279E-5 pscbe2 = 3.181440244991188E-8 lpscbe2 = -1.174751907876282E-14
+ wpscbe2 = -6.699227534670641E-14 ppscbe2 = 3.485738445798517E-20 pvag = 0
+ delta = 0.01 fprout = 0 pdits = 0
+ pditsl = 0 pditsd = 0 lambda = 0
+ vtl = 0 lc = 5E-9 xn = 3
+ alpha0 = 1E-10 alpha1 = 1E-10 beta0 = 8.93665071288678
+ lbeta0 = 8.931534583479728E-9 wbeta0 = 2.871939057542718E-6 pbeta0 = -9.913703680372806E-13
+ aigbacc = 0.43 bigbacc = 0.054 cigbacc = 0.075
+ nigbacc = 1 aigbinv = 0.35 bigbinv = 0.03
+ cigbinv = 6E-3 eigbinv = 1.1 nigbinv = 3
+ aigc = 0.43 bigc = 0.054 cigc = 0.075
+ aigsd = 0.43 bigsd = 0.054 cigsd = 0.075
+ dlcig = 0 nigc = 1 poxedge = 1
+ pigcd = 1 ntox = 1 toxref = 4.23E-9
+ agidl = 1E-10 bgidl = 7.72206191774503E8 lbgidl = 181.1931661322146
+ wbgidl = 1.770579024169947E3 pbgidl = -8.062262909721585E-4 cgidl = 300
+ egidl = 0.1 noia = 1.2E41 noib = 2E25
+ noic = 0 em = 4.1E7 af = 1
+ ef = 0.88 kf = 0 lintnoi = -6E-8
+ tnoia = 1.5 tnoib = 3.5 ntnoi = 1
+ rnoia = 0.577 rnoib = 0.37 xpart = 0
+ cgso = {5.932020000000001E-11/sw_func_tox_lv_ratio} cgdo = {5.932020000000001E-11/sw_func_tox_lv_ratio} cgbo = {0/sw_func_tox_lv_ratio}
+ ckappas = 0.6 cf = 1.2E-11 clc = 1E-7
+ cle = 0.6 dlc = -2.56E-9 dwc = 0
+ vfbcv = -0.1446893 noff = 4 voffcv = -0.1375
+ acde = 0.552 moin = 14.504 cgsl = {7.513892E-12/sw_func_tox_lv_ratio}
+ cgdl = {7.513892E-12/sw_func_tox_lv_ratio} ijthsrev = 0.1 ijthsfwd = 0.1
+ xjbvs = 1 bvs = 12.8 jss = 2.17E-5
+ jsws = 8.200000000000001E-10 cjs = {7.433E-04*sw_func_psd_nw_cj} mjs = 0.34629
+ mjsws = 0.26859 cjsws = {9.2435E-11*sw_func_psd_nw_cj} cjswgs = {2.4701E-10*sw_func_psd_nw_cj}
+ mjswgs = 0.70393 pbs = 0.6587 pbsws = 0.7418
+ pbswgs = 1.3925 xrcrg1 = 12 xrcrg2 = 1
+ rbpb = 50 rbpd = 50 rbps = 50
+ rbdb = 50 rbsb = 50 gbmin = 1E-12
+ tnom = 30 ute = -0.43771100719744 lute = 1.013292682032038E-7
+ wute = 1.180075128454327E-6 pute = -2.679382821442867E-13 kt1 = -0.525042138888159
+ lkt1 = 1.772973540392686E-8 wkt1 = 9.215076497194333E-8 pkt1 = -4.862399342741891E-14
+ kt1l = 0 kt2 = -1.826391978190144E-3 lkt2 = -6.527007591627067E-9
+ wkt2 = -1.289533344579596E-7 pkt2 = 1.552546260344322E-14 ua1 = 5.926249789932668E-9
+ lua1 = -1.50881436752443E-15 wua1 = -1.004401576172561E-14 pua1 = 3.864655445980503E-21
+ ub1 = -4.746666053748954E-18 lub1 = 1.281272423468189E-24 wub1 = 8.412609992147408E-24
+ pub1 = -3.427686384700616E-30 uc1 = -7.78091794252629E-10 luc1 = 2.249071454152068E-16
+ wuc1 = 2.264080504294589E-15 puc1 = -7.510047213808538E-22 at = 1.247866471660234E5
+ lat = -0.026600409498147 wat = -0.296619785283672 pat = 9.445444106025923E-8
+ prt = 0 njs = 1.2556 xtis = 2
+ tpb = 1.9551E-3 tpbsw = 1.4242E-4 tpbswg = 0
+ tcj = 1.2407E-3 tcjsw = 0 tcjswg = 2E-12
+ tvoff = 0 tvfbsdoff = 0 saref = 1.75E-6
+ sbref = 1.74E-6 wlod = 0 ku0 = 4.5E-8
+ kvsat = 0.4 kvth0 = 2.65E-8 tku0 = 0
+ llodku0 = 0 wlodku0 = 1 llodvth = 0
+ wlodvth = 1 lku0 = 0 wku0 = 2.5E-7
+ pku0 = 0 lkvth0 = 0 wkvth0 = 2.5E-7
+ pkvth0 = 0 stk2 = 0 lodk2 = 1
+ steta0 = 0 lodeta0 = 1

.model phighvt_model.23 pmos
+ level = 54 lmin = 1.8E-7 lmax = 2.5E-7 wmin = 3E-6
+ wmax = 5E-6 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 4.23E-9
+ toxm = 4.23E-9 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 9.999999999999999E22 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {9.364E-9+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {-1.176E-8-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = -5.722E-9 dwb = -1.7864E-8 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = -0.919198990894024 lvth0 = -3.828699263265303E-8
+ wvth0 = -2.166288595625854E-7 pvth0 = 6.320863192302371E-14 k1 = 1.154733366429159
+ lk1 = -7.320917920392118E-8 wk1 = -3.908683816802487E-6 pk1 = 8.964642092895509E-13
+ k2 = -0.211318587485936 lk2 = 2.037673631897143E-8 wk2 = 1.487775337403724E-6
+ pk2 = -3.336202138545178E-13 k3 = -13.778 k3b = 2
+ w0 = 0 lpe0 = 0 lpeb = 0
+ vbm = -3 dvtp0 = 0 dvtp1 = 0
+ dvt0 = 4.05 dvt1 = 0.3 dvt2 = 0.03
+ dvt0w = -4.254 dvt1w = 1.1472E6 dvt2w = -8.96E-3
+ vfbsdoff = 0 u0 = -0.010029902991125 lu0 = 3.783087244892618E-9
+ wu0 = 6.189141461596923E-8 pu0 = -1.551887206207604E-14 ua = -6.595232335496045E-9
+ lua = 1.180014362481962E-15 wua = 2.025610663601329E-14 pua = -4.912724620444482E-21
+ ub = 5.273967078128856E-18 lub = -8.906949194477497E-25 wub = -1.545719770426938E-23
+ pub = 3.730843367495314E-30 uc = 1.190954362693814E-10 luc = -3.384447956489881E-17
+ wuc = -5.10379507973332E-16 puc = 1.274601516527708E-22 ud = 0
+ up = 0 lp = 1 eu = 1.67
+ vsat = -6.847333610998427E3 lvsat = 0.027097069349879 wvsat = -0.061833688921336
+ pvsat = 7.77729824894334E-9 a0 = -0.499539295847909 la0 = 3.272696999364833E-7
+ wa0 = 3.95671893038869E-6 pa0 = -1.017880701657313E-12 ags = 2.292707650215772
+ lags = -2.122118609719139E-7 wags = 8.683796291147537E-6 pags = -1.767326221174347E-12
+ b0 = 0 b1 = 0 keta = -0.607430579027525
+ lketa = 1.251917603057004E-7 wketa = 1.660401490243347E-6 pketa = -3.869222117229208E-13
+ a1 = 0 a2 = 1.873052142483929 la2 = -2.935012220122043E-7
+ wa2 = -2.010479304916713E-6 pa2 = 5.499062994808193E-13 rdsw = 531.92
+ rdswmin = 0 rdw = 0 rdwmin = 0
+ rsw = 0 rswmin = 0 prwb = -0.32348
+ prwg = 0.02 wr = 1 voff = -0.230630790650497
+ lvoff = -1.47116040874913E-9 wvoff = 2.238343452342099E-7 pvoff = -5.769797531544286E-14
+ voffl = 0 minv = 0 nfactor = -3.503006302542612
+ lnfactor = 1.306660659024347E-6 wnfactor = 1.377870161602878E-5 pnfactor = -3.368676713572764E-12
+ eta0 = 0.49 etab = -6.25E-4 dsub = -1.19293434794185
+ ldsub = 5.790918682747153E-7 wdsub = 5.509379574455651E-6 pdsub = -1.782711466131895E-12
+ cit = 1E-5 cdsc = 0 cdscb = 0
+ cdscd = 0 pclm = 0.944175432949062 lpclm = -8.415408679106355E-8
+ wpclm = -1.744064609789881E-6 ppclm = 4.78733539366862E-13 pdiblc1 = -0.148186770992116
+ lpdiblc1 = 1.055673618070346E-7 wpdiblc1 = 8.364275731044141E-7 ppdiblc1 = -1.150061114156437E-13
+ pdiblc2 = 0.01386804803236 lpdiblc2 = -1.250285494427E-9 wpdiblc2 = -3.359363352957192E-8
+ ppdiblc2 = 8.144320473703376E-15 pdiblcb = -0.312971457420331 lpdiblcb = 7.8765953033609E-8
+ wpdiblcb = 2.588762559444871E-6 ppdiblcb = -7.080783352593612E-13 drout = 1.693827718856524
+ ldrout = -3.394200796463248E-7 wdrout = -5.875143031673982E-6 pdrout = 1.595152155163649E-12
+ pscbe1 = 7.9985266E8 pscbe2 = -2.778975791361339E-8 lpscbe2 = 4.555410863868612E-15
+ wpscbe2 = 1.085471164763795E-13 ppscbe2 = -1.315614999346528E-20 pvag = 0
+ delta = 0.01 fprout = 0 pdits = 0
+ pditsl = 0 pditsd = 0 lambda = 0
+ vtl = 0 lc = 5E-9 xn = 3
+ alpha0 = 1E-10 alpha1 = 1E-10 beta0 = 7.743796530837235
+ lbeta0 = 3.352010104576712E-7 wbeta0 = 9.1161688170467E-7 pbeta0 = -4.551830465020577E-13
+ aigbacc = 0.43 bigbacc = 0.054 cigbacc = 0.075
+ nigbacc = 1 aigbinv = 0.35 bigbinv = 0.03
+ cigbinv = 6E-3 eigbinv = 1.1 nigbinv = 3
+ aigc = 0.43 bigc = 0.054 cigc = 0.075
+ aigsd = 0.43 bigsd = 0.054 cigsd = 0.075
+ dlcig = 0 nigc = 1 poxedge = 1
+ pigcd = 1 ntox = 1 toxref = 4.23E-9
+ agidl = 1.055845634531155E-9 lagidl = -2.614428979569613E-16 wagidl = -4.761327095612274E-15
+ pagidl = 1.302318187191869E-21 bgidl = 2.300401376376079E9 lbgidl = -236.7987807600084
+ wbgidl = -3.412607654544003E3 pbgidl = 6.11478929389681E-4 cgidl = 300
+ egidl = 0.1 noia = 1.2E41 noib = 2E25
+ noic = 0 em = 4.1E7 af = 1
+ ef = 0.88 kf = 0 lintnoi = -6E-8
+ tnoia = 1.5 tnoib = 3.5 ntnoi = 1
+ rnoia = 0.577 rnoib = 0.37 xpart = 0
+ cgso = {5.932020000000001E-11/sw_func_tox_lv_ratio} cgdo = {5.932020000000001E-11/sw_func_tox_lv_ratio} cgbo = {0/sw_func_tox_lv_ratio}
+ ckappas = 0.6 cf = 1.2E-11 clc = 1E-7
+ cle = 0.6 dlc = -2.56E-9 dwc = 0
+ vfbcv = -0.1446893 noff = 4 voffcv = -0.1375
+ acde = 0.552 moin = 14.504 cgsl = {7.513892E-12/sw_func_tox_lv_ratio}
+ cgdl = {7.513892E-12/sw_func_tox_lv_ratio} ijthsrev = 0.1 ijthsfwd = 0.1
+ xjbvs = 1 bvs = 12.8 jss = 2.17E-5
+ jsws = 8.200000000000001E-10 cjs = {7.433E-04*sw_func_psd_nw_cj} mjs = 0.34629
+ mjsws = 0.26859 cjsws = {9.2435E-11*sw_func_psd_nw_cj} cjswgs = {2.4701E-10*sw_func_psd_nw_cj}
+ mjswgs = 0.70393 pbs = 0.6587 pbsws = 0.7418
+ pbswgs = 1.3925 xrcrg1 = 12 xrcrg2 = 1
+ rbpb = 50 rbpd = 50 rbps = 50
+ rbdb = 50 rbsb = 50 gbmin = 1E-12
+ tnom = 30 ute = 2.574251680333716 lute = -7.22502766090318E-7
+ wute = -7.50118774769186E-6 pute = 2.106560739739218E-12 kt1 = -0.50253202020399
+ lkt1 = 1.157276774143281E-8 wkt1 = 2.740216950838991E-7 pkt1 = -9.836933023164116E-14
+ kt1l = 0 kt2 = 0.072574133936601 lkt2 = -2.687703943984066E-8
+ wkt2 = -3.747843083368422E-7 pkt2 = 8.276515057879517E-14 ua1 = 2.565980705339542E-9
+ lua1 = -5.89713567506518E-16 wua1 = 5.691965406192268E-15 pua1 = -4.394501230683954E-22
+ ub1 = -2.786617815618363E-18 lub1 = 7.451600293747095E-25 wub1 = -4.446637674244336E-24
+ pub1 = 8.95750370108527E-32 uc1 = 1.265632041661894E-10 luc1 = -2.253408975230837E-17
+ wuc1 = -1.516968849663239E-15 puc1 = 2.831878979136912E-22 at = -5.259389146112648E4
+ lat = 0.021916715427151 wat = 0.582322481228497 pat = -1.459538476761494E-7
+ prt = 0 njs = 1.2556 xtis = 2
+ tpb = 1.9551E-3 tpbsw = 1.4242E-4 tpbswg = 0
+ tcj = 1.2407E-3 tcjsw = 0 tcjswg = 2E-12
+ tvoff = 0 tvfbsdoff = 0 saref = 1.25E-6
+ sbref = 1.24E-6 wlod = 0 ku0 = 4.5E-8
+ kvsat = 0.4 kvth0 = 2.65E-8 tku0 = 0
+ llodku0 = 0 wlodku0 = 1 llodvth = 0
+ wlodvth = 1 lku0 = 0 wku0 = 2.5E-7
+ pku0 = 0 lkvth0 = 0 wkvth0 = 2.5E-7
+ pkvth0 = 0 stk2 = 0 lodk2 = 1
+ steta0 = 0 lodeta0 = 1

.model phighvt_model.24 pmos
+ level = 54 lmin = 1.5E-7 lmax = 1.8E-7 wmin = 3E-6
+ wmax = 5E-6 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 4.23E-9
+ toxm = 4.23E-9 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 9.999999999999999E22 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {9.364E-9+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {-1.176E-8-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = -5.722E-9 dwb = -1.7864E-8 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = -1.119359313980131 lvth0 = 2.449636321831469E-9
+ wvth0 = 6.373442141615427E-7 pvth0 = -1.105919680413109E-13 k1 = 0.467497098151378
+ lk1 = 6.665714611597288E-8 wk1 = 3.365629296463615E-6 pk1 = -5.840039955223664E-13
+ k2 = -0.208446589538877 lk2 = 1.979222729678596E-8 wk2 = -1.027605906203728E-6
+ pk2 = 1.783101768444709E-13 k3 = -13.778 k3b = 2
+ w0 = 0 lpe0 = 0 lpeb = 0
+ vbm = -3 dvtp0 = 0 dvtp1 = 0
+ dvt0 = 4.05 dvt1 = 0.3 dvt2 = 0.03
+ dvt0w = -4.254 dvt1w = 1.1472E6 dvt2w = -8.96E-3
+ vfbsdoff = 0 u0 = 0.046121234031293 lu0 = -7.644792161910027E-9
+ wu0 = -9.742437864779909E-8 pu0 = 1.69050781829661E-14 ua = 9.917233190726889E-9
+ lua = -2.18060262141493E-15 wua = -2.63400599294352E-14 pua = 4.570527198955596E-21
+ ub = -7.000524153752133E-18 lub = 1.607409536064669E-24 wub = 1.864086189088853E-23
+ pub = -3.208793721311225E-30 uc = -3.73754388322476E-10 luc = 6.646031673603602E-17
+ wuc = 7.862571396679387E-16 puc = -1.364313388751807E-22 ud = 0
+ up = 0 lp = 1 eu = 1.67
+ vsat = 3.840359831549436E5 lvsat = -0.052455503278326 wvsat = -0.117288747351314
+ pvsat = 1.906351174061252E-8 a0 = 0.774149454850561 la0 = 6.804856539433068E-8
+ wa0 = -7.086975498153548E-6 pa0 = 1.229731988439604E-12 ags = 1.25
+ b0 = 0 b1 = 0 keta = 0.378072655192662
+ lketa = -7.537785792279194E-8 wketa = -2.118015585694881E-6 pketa = 3.820612315720276E-13
+ a1 = 0 a2 = 0.306175092737501 la2 = 2.538959515218884E-8
+ wa2 = 4.691118378138986E-6 pa2 = -8.140028609746767E-13 rdsw = 531.92
+ rdswmin = 0 rdw = 0 rdwmin = 0
+ rsw = 0 rswmin = 0 prwb = -0.32348
+ prwg = 0.02 wr = 1 voff = -0.10275322558461
+ lvoff = -2.749680245095855E-8 wvoff = -4.047736457792144E-7 pvoff = 7.023632301560928E-14
+ voffl = 0 minv = 0 nfactor = 8.670871190762481
+ lnfactor = -1.170966888413106E-6 wnfactor = -1.881451202261953E-5 pnfactor = 3.264694126164941E-12
+ eta0 = 0.49 etab = -4.203849999999993E-3 letab = 7.283675519999987E-10
+ dsub = 7.380402828426323 ldsub = -1.165753713859736E-6 wdsub = -2.204808450462265E-5
+ pdsub = 3.825783623242121E-12 cit = 1E-5 cdsc = 0
+ cdscb = 0 cdscd = 0 pclm = -1.181247596122344
+ lpclm = 3.484120080855491E-7 wpclm = 4.126050332747507E-6 ppclm = -7.159522537383473E-13
+ pdiblc1 = 1.427562604623973 lpdiblc1 = -2.151291511183517E-7 wpdiblc1 = 1.840787608752219E-6
+ ppdiblc1 = -3.194134658706849E-13 pdiblc2 = -0.156685822621636 lpdiblc2 = 3.346083826107429E-8
+ wpdiblc2 = 4.357813925882982E-8 ppdiblc2 = -7.56167872419215E-15 pdiblcb = 1.803733400647437
+ lpdiblcb = -3.520258196803432E-7 wpdiblcb = -6.04044597203802E-6 ppdiblcb = 1.048138185068037E-12
+ drout = -5.596110681354823 ldrout = 1.144228183564689E-6 wdrout = 1.331476817857864E-5
+ pdrout = -2.310378574346966E-12 pscbe1 = 8E8 pscbe2 = -9.057100651353274E-8
+ lpscbe2 = 1.73326505789242E-14 wpscbe2 = 2.978453050602488E-13 ppscbe2 = -5.168211733405436E-20
+ pvag = 0 delta = 0.01 fprout = 0
+ pdits = 0 pditsl = 0 pditsd = 0
+ lambda = 0 vtl = 0 lc = 5E-9
+ xn = 3 alpha0 = 1E-10 alpha1 = 1E-10
+ beta0 = 11.158402012455518 lbeta0 = -3.597394971612812E-7 wbeta0 = -8.988359291250759E-6
+ pbeta0 = 1.559660104217831E-12 aigbacc = 0.43 bigbacc = 0.054
+ cigbacc = 0.075 nigbacc = 1 aigbinv = 0.35
+ bigbinv = 0.03 cigbinv = 6E-3 eigbinv = 1.1
+ nigbinv = 3 aigc = 0.43 bigc = 0.054
+ cigc = 0.075 aigsd = 0.43 bigsd = 0.054
+ cigsd = 0.075 dlcig = 0 nigc = 1
+ poxedge = 1 pigcd = 1 ntox = 1
+ toxref = 4.23E-9 agidl = -1.420090277372701E-9 lagidl = 2.424595788337114E-16
+ wagidl = 6.814990890470367E-15 pagidl = -1.05369404933567E-21 bgidl = 1.928630245335038E9
+ lbgidl = -161.13592017053585 wbgidl = -2.768499348770481E3 pbgidl = 4.803900069986538E-4
+ cgidl = 300 egidl = 0.1 noia = 1.2E41
+ noib = 2E25 noic = 0 em = 4.1E7
+ af = 1 ef = 0.88 kf = 0
+ lintnoi = -6E-8 tnoia = 1.5 tnoib = 3.5
+ ntnoi = 1 rnoia = 0.577 rnoib = 0.37
+ xpart = 0 cgso = {5.932020000000001E-11/sw_func_tox_lv_ratio} cgdo = {5.932020000000001E-11/sw_func_tox_lv_ratio}
+ cgbo = {0/sw_func_tox_lv_ratio} ckappas = 0.6 cf = 1.2E-11
+ clc = 1E-7 cle = 0.6 dlc = -2.56E-9
+ dwc = 0 vfbcv = -0.1446893 noff = 4
+ voffcv = -0.1375 acde = 0.552 moin = 14.504
+ cgsl = {7.513892E-12/sw_func_tox_lv_ratio} cgdl = {7.513892E-12/sw_func_tox_lv_ratio} ijthsrev = 0.1
+ ijthsfwd = 0.1 xjbvs = 1 bvs = 12.8
+ jss = 2.17E-5 jsws = 8.200000000000001E-10 cjs = {7.433E-04*sw_func_psd_nw_cj}
+ mjs = 0.34629 mjsws = 0.26859 cjsws = {9.2435E-11*sw_func_psd_nw_cj}
+ cjswgs = {2.4701E-10*sw_func_psd_nw_cj} mjswgs = 0.70393 pbs = 0.6587
+ pbsws = 0.7418 pbswgs = 1.3925 xrcrg1 = 12
+ xrcrg2 = 1 rbpb = 50 rbpd = 50
+ rbps = 50 rbdb = 50 rbsb = 50
+ gbmin = 1E-12 tnom = 30 ute = -6.51568730815999
+ lute = 1.127481616847922E-6 wute = 2.147801981061147E-5 pute = -3.791287582526676E-12
+ kt1 = 0.251561393410558 lkt1 = -1.419003237974E-7 wkt1 = -9.90537261676365E-7
+ pkt1 = 1.589937086482079E-13 kt1l = 0 kt2 = -0.158704318035456
+ lkt2 = 2.019275110551229E-8 wkt2 = 2.163016048693676E-7 pkt2 = -3.753265447693267E-14
+ ua1 = -3.946126531860473E-9 lua1 = 7.356304974084295E-16 wua1 = 2.396595587999512E-14
+ pua1 = -4.158572664296753E-21 ub1 = 5.618596368668663E-18 lub1 = -9.654691614113867E-25
+ wub1 = -2.71801554150451E-23 pub1 = 4.716300567618626E-30 uc1 = 4.448780919864824E-10
+ luc1 = -8.731753572149442E-17 wuc1 = -8.515200789923736E-16 puc1 = 1.477557641067567E-22
+ at = -8.86553090072573E4 lat = 0.029255935126139 wat = -0.485175309955023
+ pat = 7.130330278552072E-8 prt = 0 njs = 1.2556
+ xtis = 2 tpb = 1.9551E-3 tpbsw = 1.4242E-4
+ tpbswg = 0 tcj = 1.2407E-3 tcjsw = 0
+ tcjswg = 2E-12 tvoff = 0 tvfbsdoff = 0
+ saref = 1.1E-6 sbref = 1.1E-6 wlod = 0
+ ku0 = 4.5E-8 kvsat = 0.4 kvth0 = 2.65E-8
+ tku0 = 0 llodku0 = 0 wlodku0 = 1
+ llodvth = 0 wlodvth = 1 lku0 = 0
+ wku0 = 2.5E-7 pku0 = 0 lkvth0 = 0
+ wkvth0 = 2.5E-7 pkvth0 = 0 stk2 = 0
+ lodk2 = 1 steta0 = 0 lodeta0 = 1

.model phighvt_model.25 pmos
+ level = 54 lmin = 8E-6 lmax = 2.02E-5 wmin = 1E-6
+ wmax = 3E-6 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 4.23E-9
+ toxm = 4.23E-9 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 9.999999999999999E22 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {9.364E-9+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {-1.176E-8-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = -5.722E-9 dwb = -1.7864E-8 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = -1.0761835273908 wvth0 = -1.177445210457481E-8
+ k1 = 0.50470237751996 wk1 = -5.611373269208613E-8 k2 = 9.216488098376002E-3
+ wk2 = 1.154821915065038E-8 k3 = -13.778 k3b = 2
+ w0 = 0 lpe0 = 0 lpeb = 0
+ vbm = -3 dvtp0 = 0 dvtp1 = 0
+ dvt0 = 4.05 dvt1 = 0.3 dvt2 = 0.03
+ dvt0w = -4.254 dvt1w = 1.1472E6 dvt2w = -8.96E-3
+ vfbsdoff = 0 u0 = 7.9909699790936E-3 wu0 = 1.008482693074864E-9
+ ua = -6.521572587540017E-11 wua = -6.491107549696743E-16 ub = -1.884280847276399E-19
+ wub = 1.15171815620878E-24 uc = -1.27564678295916E-10 wuc = 5.474297595254208E-17
+ ud = 0 up = 0 lp = 1
+ eu = 1.67 vsat = 1.6031E5 a0 = 1.831927806302
+ wa0 = -5.657718069695759E-7 ags = 0.5354464690062 wags = -2.869057488546518E-7
+ b0 = 0 b1 = 0 keta = -0.0456438813829
+ wketa = 4.295388787796104E-8 a1 = 0 a2 = 0.8
+ rdsw = 531.92 rdswmin = 0 rdw = 0
+ rdwmin = 0 rsw = 0 rswmin = 0
+ prwb = -0.32348 prwg = 0.02 wr = 1
+ voff = -0.1709520165572 wvoff = -4.030859646712324E-8 voffl = 0
+ minv = 0 nfactor = 2.848616973416 wnfactor = -1.014550930649065E-6
+ eta0 = 0.08 etab = -0.07 dsub = 0.56
+ cit = 1E-5 cdsc = 0 cdscb = 0
+ cdscd = 0 pclm = 0.02049648869966 wpclm = 1.182064697632672E-7
+ pdiblc1 = 0.39 pdiblc2 = 2.7113785151308E-4 wpdiblc2 = 4.725822485149697E-11
+ pdiblcb = 0.073826071761906 wpdiblcb = -2.246579085321094E-7 drout = 0.56
+ pscbe1 = 7.855045276106E8 wpscbe1 = 14.176164172491314 pscbe2 = 1.12912238292372E-8
+ wpscbe2 = -5.755907056681644E-15 pvag = 0 delta = 0.01
+ fprout = 0 pdits = 0 pditsl = 0
+ pditsd = 0 lambda = 0 vtl = 0
+ lc = 5E-9 xn = 3 alpha0 = 1E-10
+ alpha1 = 1E-10 beta0 = 1.391406060205201 wbeta0 = 4.795656072079922E-6
+ aigbacc = 0.43 bigbacc = 0.054 cigbacc = 0.075
+ nigbacc = 1 aigbinv = 0.35 bigbinv = 0.03
+ cigbinv = 6E-3 eigbinv = 1.1 nigbinv = 3
+ aigc = 0.43 bigc = 0.054 cigc = 0.075
+ aigsd = 0.43 bigsd = 0.054 cigsd = 0.075
+ dlcig = 0 nigc = 1 poxedge = 1
+ pigcd = 1 ntox = 1 toxref = 4.23E-9
+ agidl = -8.497305123999656E-13 wagidl = 4.375957564719237E-16 bgidl = 1E9
+ cgidl = 300 egidl = -0.2853698744774 wegidl = 1.148892416422987E-6
+ noia = 1.2E41 noib = 2E25 noic = 0
+ em = 4.1E7 af = 1 ef = 0.88
+ kf = 0 lintnoi = -6E-8 tnoia = 1.5
+ tnoib = 3.5 ntnoi = 1 rnoia = 0.577
+ rnoib = 0.37 xpart = 0 cgso = {5.932020000000001E-11/sw_func_tox_lv_ratio}
+ cgdo = {5.932020000000001E-11/sw_func_tox_lv_ratio} cgbo = {0/sw_func_tox_lv_ratio} ckappas = 0.6
+ cf = 1.2E-11 clc = 1E-7 cle = 0.6
+ dlc = -2.56E-9 dwc = 0 vfbcv = -0.1446893
+ noff = 4 voffcv = -0.1375 acde = 0.552
+ moin = 14.504 cgsl = {7.513892E-12/sw_func_tox_lv_ratio} cgdl = {7.513892E-12/sw_func_tox_lv_ratio}
+ ijthsrev = 0.1 ijthsfwd = 0.1 xjbvs = 1
+ bvs = 12.8 jss = 2.17E-5 jsws = 8.200000000000001E-10
+ cjs = {7.433E-04*sw_func_psd_nw_cj} mjs = 0.34629 mjsws = 0.26859
+ cjsws = {9.2435E-11*sw_func_psd_nw_cj} cjswgs = {2.4701E-10*sw_func_psd_nw_cj} mjswgs = 0.70393
+ pbs = 0.6587 pbsws = 0.7418 pbswgs = 1.3925
+ xrcrg1 = 12 xrcrg2 = 1 rbpb = 50
+ rbpd = 50 rbps = 50 rbdb = 50
+ rbsb = 50 gbmin = 1E-12 tnom = 30
+ ute = -0.42655326278768 wute = 2.887757331775523E-7 kt1 = -0.462785957766
+ wkt1 = 2.160217100095837E-8 kt1l = 0 kt2 = -0.030897081927808
+ wkt2 = -2.105946115891999E-8 ua1 = 2.8309542679452E-9 wua1 = -9.893478371055224E-16
+ ub1 = -2.15422013227232E-18 wub1 = 1.411394184579764E-24 uc1 = 6.391306549818012E-10
+ wuc1 = -6.357582066789043E-16 at = 0 prt = 0
+ njs = 1.2556 xtis = 2 tpb = 1.9551E-3
+ tpbsw = 1.4242E-4 tpbswg = 0 tcj = 1.2407E-3
+ tcjsw = 0 tcjswg = 2E-12 tvoff = 0
+ tvfbsdoff = 0 saref = 3E-6 sbref = 3E-6
+ wlod = 0 ku0 = 4.5E-8 kvsat = 0.4
+ kvth0 = 2.65E-8 tku0 = 0 llodku0 = 0
+ wlodku0 = 1 llodvth = 0 wlodvth = 1
+ lku0 = 0 wku0 = 2.5E-7 pku0 = 0
+ lkvth0 = 0 wkvth0 = 2.5E-7 pkvth0 = 0
+ stk2 = 0 lodk2 = 1 steta0 = 0
+ lodeta0 = 1

.model phighvt_model.26 pmos
+ level = 54 lmin = 4E-6 lmax = 8E-6 wmin = 1E-6
+ wmax = 3E-6 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 4.23E-9
+ toxm = 4.23E-9 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 9.999999999999999E22 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {9.364E-9+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {-1.176E-8-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = -5.722E-9 dwb = -1.7864E-8 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = -1.094894426939826 lvth0 = 1.501272767495974E-7
+ wvth0 = 4.32261437287981E-9 pvth0 = -1.291551348231867E-13 k1 = 0.450206226023736
+ lk1 = 4.372509614529834E-7 wk1 = 5.364276656665435E-9 pk1 = -4.932700375698951E-13
+ k2 = 0.022658357815787 lk2 = -1.078511105150449E-7 wk2 = -3.733123301069486E-9
+ pk2 = 1.226101567882234E-13 k3 = -13.778 k3b = 2
+ w0 = 0 lpe0 = 0 lpeb = 0
+ vbm = -3 dvtp0 = 0 dvtp1 = 0
+ dvt0 = 4.05 dvt1 = 0.3 dvt2 = 0.03
+ dvt0w = -4.254 dvt1w = 1.1472E6 dvt2w = -8.96E-3
+ vfbsdoff = 0 u0 = 0.011641682507783 lu0 = -2.929156498818803E-8
+ wu0 = -3.04724457671806E-9 pu0 = 3.254120886372893E-14 ua = 9.669688893892674E-10
+ lua = -8.281753904268364E-15 wua = -1.757219053845627E-15 pua = 8.89092909819718E-21
+ ub = -8.66101985372604E-19 lub = 5.437330095302884E-24 wub = 1.878763641406163E-24
+ pub = -5.833463991390903E-30 uc = -1.778366324767365E-10 luc = 4.033580298088972E-16
+ wuc = 1.049947418656588E-16 puc = -4.031960488392105E-22 ud = 0
+ up = 0 lp = 1 eu = 1.67
+ vsat = 1.992067948535321E5 lvsat = -0.312059311073815 wvsat = 0.067318804051447
+ pvsat = -5.40163111078143E-7 a0 = 1.836036115254248 la0 = -3.296309904454598E-8
+ wa0 = -4.834942594967697E-7 pa0 = -6.601555476990101E-13 ags = 0.567879070176478
+ lags = -2.602236241417503E-7 wags = -3.559878350485355E-7 pags = 5.542815002183499E-13
+ b0 = 0 b1 = 0 keta = -0.055472811009576
+ lketa = 7.886261343822907E-8 wketa = 5.361312425000713E-8 pketa = -8.55245962158392E-14
+ a1 = 0 a2 = 0.8 rdsw = 531.92
+ rdswmin = 0 rdw = 0 rdwmin = 0
+ rsw = 0 rswmin = 0 prwb = -0.32348
+ prwg = 0.02 wr = 1 voff = -0.183949195662276
+ lvoff = 1.042831264931625E-7 wvoff = -2.136989580081267E-8 pvoff = -1.519550435701562E-13
+ voffl = 0 minv = 0 nfactor = 2.980137016766105
+ lnfactor = -1.055253698220435E-6 wnfactor = -8.143614913794493E-7 pnfactor = -1.606223969768546E-12
+ eta0 = 0.08 etab = -0.07 dsub = 0.56
+ cit = 1E-5 cdsc = 0 cdscb = 0
+ cdscd = 0 pclm = -0.887103000636486 lpclm = 7.282142654678351E-6
+ wpclm = 1.106694532891214E-6 ppclm = -7.93115374426834E-12 pdiblc1 = 0.39
+ pdiblc2 = 1.221485478409193E-3 lpdiblc2 = -7.625133191353502E-9 wpdiblc2 = -2.570104147646051E-9
+ ppdiblc2 = 2.100045934298153E-14 pdiblcb = 0.121714603232206 lpdiblcb = -3.842345900225739E-7
+ wpdiblcb = -3.641657325687243E-7 ppdiblcb = 1.11934381631426E-12 drout = 0.56
+ pscbe1 = 5.612699823317872E8 lpscbe1 = 1.799150358735459E3 wpscbe1 = 653.4708056192295
+ ppscbe1 = -5.129393341540733E-3 pscbe2 = 2.203884114376791E-8 lpscbe2 = -8.623372247548339E-14
+ wpscbe2 = -3.842154868615483E-14 ppscbe2 = 2.620934289269107E-19 pvag = 0
+ delta = 0.01 fprout = 0 pdits = 0
+ pditsl = 0 pditsd = 0 lambda = 0
+ vtl = 0 lc = 5E-9 xn = 3
+ alpha0 = 1E-10 alpha1 = 1E-10 beta0 = -2.746899343935037
+ lbeta0 = 3.320377617622728E-5 wbeta0 = 6.060802638341774E-6 pbeta0 = -1.01509287773333E-11
+ aigbacc = 0.43 bigbacc = 0.054 cigbacc = 0.075
+ nigbacc = 1 aigbinv = 0.35 bigbinv = 0.03
+ cigbinv = 6E-3 eigbinv = 1.1 nigbinv = 3
+ aigc = 0.43 bigc = 0.054 cigc = 0.075
+ aigsd = 0.43 bigsd = 0.054 cigsd = 0.075
+ dlcig = 0 nigc = 1 poxedge = 1
+ pigcd = 1 ntox = 1 toxref = 4.23E-9
+ agidl = -5.309021123512787E-11 lagidl = 4.19152541888422E-16 wagidl = 7.310792970435763E-16
+ pagidl = -2.354771057447466E-21 bgidl = 7.026774901869061E8 lbgidl = 2.385573103935555E3
+ wbgidl = 291.7542538493141 pbgidl = -2.340896090845049E-3 cgidl = 300
+ egidl = -0.673005723816727 legidl = 3.110203989891076E-6 wegidl = 2.304540320254541E-6
+ pegidl = -9.272364069350551E-12 noia = 1.2E41 noib = 2E25
+ noic = 0 em = 4.1E7 af = 1
+ ef = 0.88 kf = 0 lintnoi = -6E-8
+ tnoia = 1.5 tnoib = 3.5 ntnoi = 1
+ rnoia = 0.577 rnoib = 0.37 xpart = 0
+ cgso = {5.932020000000001E-11/sw_func_tox_lv_ratio} cgdo = {5.932020000000001E-11/sw_func_tox_lv_ratio} cgbo = {0/sw_func_tox_lv_ratio}
+ ckappas = 0.6 cf = 1.2E-11 clc = 1E-7
+ cle = 0.6 dlc = -2.56E-9 dwc = 0
+ vfbcv = -0.1446893 noff = 4 voffcv = -0.1375
+ acde = 0.552 moin = 14.504 cgsl = {7.513892E-12/sw_func_tox_lv_ratio}
+ cgdl = {7.513892E-12/sw_func_tox_lv_ratio} ijthsrev = 0.1 ijthsfwd = 0.1
+ xjbvs = 1 bvs = 12.8 jss = 2.17E-5
+ jsws = 8.200000000000001E-10 cjs = {7.433E-04*sw_func_psd_nw_cj} mjs = 0.34629
+ mjsws = 0.26859 cjsws = {9.2435E-11*sw_func_psd_nw_cj} cjswgs = {2.4701E-10*sw_func_psd_nw_cj}
+ mjswgs = 0.70393 pbs = 0.6587 pbsws = 0.7418
+ pbswgs = 1.3925 xrcrg1 = 12 xrcrg2 = 1
+ rbpb = 50 rbpd = 50 rbps = 50
+ rbdb = 50 rbsb = 50 gbmin = 1E-12
+ tnom = 30 ute = 0.328260532139455 lute = -6.056263579873764E-6
+ wute = -4.837499207226424E-7 pute = 6.19837503458129E-12 kt1 = -0.561884150513443
+ lkt1 = 7.951163314729662E-7 wkt1 = 1.528564353945541E-7 pkt1 = -1.053121215447303E-12
+ kt1l = 0 kt2 = -0.022961749858592 lkt2 = -6.366929556399989E-8
+ wkt2 = -2.495474008259477E-8 pkt2 = 3.125384834968313E-14 ua1 = 7.699060729150728E-9
+ lua1 = -3.905934955361178E-14 wua1 = -6.995226259379061E-15 pua1 = 4.818828563868018E-20
+ ub1 = -6.734394385632452E-18 lub1 = 3.67491197253201E-23 wub1 = 7.416765619352955E-24
+ pub1 = -4.81842178143314E-29 uc1 = 1.188188442729139E-9 luc1 = -4.405376141146521E-15
+ wuc1 = -1.17736641725454E-15 puc1 = 4.345604309717823E-21 at = -2.242570178615651E5
+ lat = 1.799330667952625 wat = 0.130556122978206 pat = -1.047519663838098E-6
+ prt = 0 njs = 1.2556 xtis = 2
+ tpb = 1.9551E-3 tpbsw = 1.4242E-4 tpbswg = 0
+ tcj = 1.2407E-3 tcjsw = 0 tcjswg = 2E-12
+ tvoff = 0 tvfbsdoff = 0 saref = 3E-6
+ sbref = 3E-6 wlod = 0 ku0 = 4.5E-8
+ kvsat = 0.4 kvth0 = 2.65E-8 tku0 = 0
+ llodku0 = 0 wlodku0 = 1 llodvth = 0
+ wlodvth = 1 lku0 = 0 wku0 = 2.5E-7
+ pku0 = 0 lkvth0 = 0 wkvth0 = 2.5E-7
+ pkvth0 = 0 stk2 = 0 lodk2 = 1
+ steta0 = 0 lodeta0 = 1

.model phighvt_model.27 pmos
+ level = 54 lmin = 2E-6 lmax = 4E-6 wmin = 1E-6
+ wmax = 3E-6 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 4.23E-9
+ toxm = 4.23E-9 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 9.999999999999999E22 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {9.364E-9+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {-1.176E-8-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = -5.722E-9 dwb = -1.7864E-8 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = -1.022821560625115 lvth0 = -1.398593423249678E-7
+ wvth0 = -6.134546165892955E-8 pvth0 = 1.350616824523189E-13 k1 = 0.67581002810476
+ lk1 = -4.704704482960608E-7 wk1 = -2.286390968010963E-7 pk1 = 4.482472156048784E-13
+ k2 = -0.030131037369593 lk2 = 1.04548076801235E-7 wk2 = 5.10894305385072E-8
+ pk2 = -9.79694850363902E-14 k3 = -13.778 k3b = 2
+ w0 = 0 lpe0 = 0 lpeb = 0
+ vbm = -3 dvtp0 = 0 dvtp1 = 0
+ dvt0 = 4.05 dvt1 = 0.3 dvt2 = 0.03
+ dvt0w = -4.254 dvt1w = 1.1472E6 dvt2w = -8.96E-3
+ vfbsdoff = 0 u0 = 9.442994008218046E-4 lu0 = 1.374956989033151E-8
+ wu0 = 7.545741471658164E-9 pu0 = -1.007988236163378E-14 ua = -1.77272037527114E-9
+ lua = 2.741440645878079E-15 wua = 9.333433709404682E-16 pua = -1.934602629178167E-21
+ ub = 7.934833502153631E-19 lub = -1.240044694142015E-24 wub = 2.139377294498202E-25
+ pub = 8.649963618836814E-31 uc = -6.246907621636202E-11 luc = -6.08256401558449E-17
+ wuc = -1.288875746859416E-17 puc = 7.11105684021431E-23 ud = 0
+ up = 0 lp = 1 eu = 1.67
+ vsat = 1.906601751976342E5 lvsat = -0.277671815955917 wvsat = -0.134652278300533
+ pvsat = 2.724715781866944E-7 a0 = 2.481176407449544 la0 = -2.628697967498163E-6
+ wa0 = -1.281204388328521E-6 pa0 = 2.549447109858117E-12 ags = 0.701108656956467
+ lags = -7.962755311427715E-7 wags = -5.286984787477205E-7 pags = 1.249186229354894E-12
+ b0 = 0 b1 = 0 keta = -0.065035975779155
+ lketa = 1.173401981519245E-7 wketa = 7.027312810931031E-8 pketa = -1.525564549438228E-13
+ a1 = 0 a2 = 0.8 rdsw = 531.92
+ rdswmin = 0 rdw = 0 rdwmin = 0
+ rsw = 0 rswmin = 0 prwb = -0.32348
+ prwg = 0.02 wr = 1 voff = -0.097149071708622
+ lvoff = -2.449589082368454E-7 wvoff = -1.340777282957072E-7 pvoff = 3.015271746297018E-13
+ voffl = 0 minv = 0 nfactor = 4.36778726734016
+ lnfactor = -6.638492234410159E-6 wnfactor = -3.512580713391822E-6 pnfactor = 9.250115034382675E-12
+ eta0 = 0.04053573259088 leta0 = 1.587852692059424E-7 weta0 = 1.17653715427322E-7
+ peta0 = -4.733820770961385E-13 etab = -0.035499171467854 letab = -1.388147736156609E-7
+ wetab = -1.028563540796886E-7 petab = 4.138445977667086E-13 dsub = 0.41172306246523
+ ldsub = 5.965952237098985E-7 wdsub = 4.420538821181594E-7 pdsub = -1.778612635780056E-12
+ cit = 1E-5 cdsc = 0 cdscb = 0
+ cdscd = 0 pclm = 1.672282372300624 lpclm = -3.015595581041568E-6
+ wpclm = -2.18652402701583E-6 ppclm = 5.319176995888846E-12 pdiblc1 = 0.39
+ pdiblc2 = -1.466032105569874E-3 lpdiblc2 = 3.188147558137948E-9 wpdiblc2 = 5.011613947436506E-9
+ ppdiblc2 = -9.504735046945038E-15 pdiblcb = 0.078037275187135 lpdiblcb = -2.084979870866707E-7
+ wpdiblcb = -1.729421459953266E-7 ppdiblcb = 3.499518912644633E-13 drout = 0.56
+ pscbe1 = 1.215455802710456E9 lpscbe1 = -832.9793732745205 wpscbe1 = -1.238586751858206E3
+ ppscbe1 = 2.483338082120877E-3 pscbe2 = 2.275258131848406E-9 lpscbe2 = -6.714550955365074E-15
+ wpscbe2 = 4.343192181052928E-14 ppscbe2 = -6.724564668590779E-20 pvag = 0
+ delta = 0.01 fprout = 0 pdits = 0
+ pditsl = 0 pditsd = 0 lambda = 0
+ vtl = 0 lc = 5E-9 xn = 3
+ alpha0 = 1E-10 alpha1 = 1E-10 beta0 = 2.638195535547811
+ lbeta0 = 1.153673922673046E-5 wbeta0 = 8.669926110399809E-6 pbeta0 = -2.064878924962824E-11
+ aigbacc = 0.43 bigbacc = 0.054 cigbacc = 0.075
+ nigbacc = 1 aigbinv = 0.35 bigbinv = 0.03
+ cigbinv = 6E-3 eigbinv = 1.1 nigbinv = 3
+ aigc = 0.43 bigc = 0.054 cigc = 0.075
+ aigsd = 0.43 bigsd = 0.054 cigsd = 0.075
+ dlcig = 0 nigc = 1 poxedge = 1
+ pigcd = 1 ntox = 1 toxref = 4.23E-9
+ agidl = 1.663622350191098E-11 lagidl = 1.386068371952513E-16 wagidl = 2.485300926880108E-16
+ pagidl = -4.132246827387612E-22 bgidl = 1.211745833510753E9 lbgidl = 337.3264432051885
+ wbgidl = -207.78025754076404 pbgidl = -3.310089935768418E-4 cgidl = 300
+ egidl = 0.1 noia = 1.2E41 noib = 2E25
+ noic = 0 em = 4.1E7 af = 1
+ ef = 0.88 kf = 0 lintnoi = -6E-8
+ tnoia = 1.5 tnoib = 3.5 ntnoi = 1
+ rnoia = 0.577 rnoib = 0.37 xpart = 0
+ cgso = {5.932020000000001E-11/sw_func_tox_lv_ratio} cgdo = {5.932020000000001E-11/sw_func_tox_lv_ratio} cgbo = {0/sw_func_tox_lv_ratio}
+ ckappas = 0.6 cf = 1.2E-11 clc = 1E-7
+ cle = 0.6 dlc = -2.56E-9 dwc = 0
+ vfbcv = -0.1446893 noff = 4 voffcv = -0.1375
+ acde = 0.552 moin = 14.504 cgsl = {7.513892E-12/sw_func_tox_lv_ratio}
+ cgdl = {7.513892E-12/sw_func_tox_lv_ratio} ijthsrev = 0.1 ijthsfwd = 0.1
+ xjbvs = 1 bvs = 12.8 jss = 2.17E-5
+ jsws = 8.200000000000001E-10 cjs = {7.433E-04*sw_func_psd_nw_cj} mjs = 0.34629
+ mjsws = 0.26859 cjsws = {9.2435E-11*sw_func_psd_nw_cj} cjswgs = {2.4701E-10*sw_func_psd_nw_cj}
+ mjswgs = 0.70393 pbs = 0.6587 pbsws = 0.7418
+ pbswgs = 1.3925 xrcrg1 = 12 xrcrg2 = 1
+ rbpb = 50 rbpd = 50 rbps = 50
+ rbdb = 50 rbsb = 50 gbmin = 1E-12
+ tnom = 30 ute = -2.401328764697562 lute = 4.926293547735906E-6
+ wute = 2.226105069515402E-6 pute = -4.704780715741287E-12 kt1 = -0.27422403697283
+ lkt1 = -3.622898885599641E-7 wkt1 = -2.035061655491208E-7 pkt1 = 3.807108367015916E-13
+ kt1l = 0 kt2 = -0.030191896397676 lkt2 = -3.457865636106439E-8
+ wkt2 = -2.953081782765817E-8 pkt2 = 4.966578867850059E-14 ua1 = -6.588130010284021E-9
+ lua1 = 1.842544813031872E-14 wua1 = 9.72617584683171E-15 pua1 = -1.909061016370098E-20
+ ub1 = 6.179823212837813E-18 lub1 = -1.521149306647698E-23 wub1 = -8.853179568466248E-24
+ pub1 = 1.727823204776292E-29 uc1 = 1.292801162682473E-10 luc1 = -1.44837311464594E-16
+ wuc1 = -1.090144855838986E-16 puc1 = 4.706894560236492E-23 at = 3.61607107216717E5
+ lat = -0.557905356582345 wat = -0.254455659203622 pat = 5.01582942006131E-7
+ prt = 0 njs = 1.2556 xtis = 2
+ tpb = 1.9551E-3 tpbsw = 1.4242E-4 tpbswg = 0
+ tcj = 1.2407E-3 tcjsw = 0 tcjswg = 2E-12
+ tvoff = 0 tvfbsdoff = 0 saref = 3E-6
+ sbref = 3E-6 wlod = 0 ku0 = 4.5E-8
+ kvsat = 0.4 kvth0 = 2.65E-8 tku0 = 0
+ llodku0 = 0 wlodku0 = 1 llodvth = 0
+ wlodvth = 1 lku0 = 0 wku0 = 2.5E-7
+ pku0 = 0 lkvth0 = 0 wkvth0 = 2.5E-7
+ pkvth0 = 0 stk2 = 0 lodk2 = 1
+ steta0 = 0 lodeta0 = 1

.model phighvt_model.28 pmos
+ level = 54 lmin = 1E-6 lmax = 2E-6 wmin = 1E-6
+ wmax = 3E-6 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 4.23E-9
+ toxm = 4.23E-9 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 9.999999999999999E22 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {9.364E-9+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {-1.176E-8-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = -5.722E-9 dwb = -1.7864E-8 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = -1.101885177433208 lvth0 = 2.012746755854489E-8
+ wvth0 = 2.845703962693229E-10 pvth0 = 1.035207998798289E-14 k1 = 0.470245475147659
+ lk1 = -5.450646409630738E-8 wk1 = -1.140363697922904E-7 pk1 = 2.163463054480197E-13
+ k2 = 0.011788787318025 lk2 = 1.972247314934776E-8 wk2 = 4.316489167686377E-8
+ pk2 = -8.193402215907747E-14 k3 = -13.778 k3b = 2
+ w0 = 0 lpe0 = 0 lpeb = 0
+ vbm = -3 dvtp0 = 0 dvtp1 = 0
+ dvt0 = 4.05 dvt1 = 0.3 dvt2 = 0.03
+ dvt0w = -4.254 dvt1w = 1.1472E6 dvt2w = -8.96E-3
+ vfbsdoff = 0 u0 = 6.77939330170097E-3 lu0 = 1.942140680024502E-9
+ wu0 = 5.616834269953448E-9 pu0 = -6.176700060840256E-15 ua = -9.28301277414768E-11
+ lua = -6.578508678031459E-16 wua = 1.16928729419608E-16 pua = -2.825712737678763E-22
+ ub = -5.130236428056583E-19 lub = 1.403698336375883E-24 wub = 1.089915319994515E-24
+ pub = -9.075618121353201E-31 uc = -1.460859249230217E-10 luc = 1.083747255390551E-16
+ wuc = 6.966459998285628E-17 puc = -9.593780146801588E-23 ud = 0
+ up = 0 lp = 1 eu = 1.67
+ vsat = 3.025205815129408E4 lvsat = 0.046917217049693 wvsat = 0.028836077022415
+ pvsat = -5.835037857639692E-8 a0 = 1.043638313826983 la0 = 2.801891157089617E-7
+ wa0 = 3.174724437495071E-7 pa0 = -6.855074333884139E-13 ags = 0.047426524807314
+ lags = 5.264633369036827E-7 wags = 1.256917680641176E-7 pags = -7.498552287379614E-14
+ b0 = 0 b1 = 0 keta = 1.699443239898175E-3
+ lketa = -1.770025694150986E-8 wketa = -1.226470885344472E-8 pketa = 1.446050890705132E-14
+ a1 = 0 a2 = 0.900435151744 la2 = -2.032325382570188E-7
+ wa2 = -2.994245057101382E-7 pa2 = 6.058914757945789E-13 rdsw = 531.92
+ rdswmin = 0 rdw = 0 rdwmin = 0
+ rsw = 0 rswmin = 0 prwb = -0.32348
+ prwg = 0.02 wr = 1 voff = -0.231534651508023
+ lvoff = 2.697300019883838E-8 wvoff = 2.880853426711434E-8 pvoff = -2.807643539141883E-14
+ voffl = 0 minv = 0 nfactor = 0.434607456515247
+ lnfactor = 1.320375776390271E-6 wnfactor = 1.958486271921939E-6 pnfactor = -1.820698431739427E-12
+ eta0 = 0.017168265693959 leta0 = 2.060698058211999E-7 weta0 = -2.368112604921226E-7
+ peta0 = 2.438848909763758E-13 etab = 0.645184592491903 letab = -1.516191983663508E-6
+ wetab = 1.953859611805173E-7 petab = -1.896546920086232E-13 dsub = 0.705697455314829
+ ldsub = 1.732160290878182E-9 wdsub = -9.537983688035946E-7 pdsub = 1.045922311005131E-12
+ cit = 1E-5 cdsc = 0 cdscb = 0
+ cdscd = 0 pclm = -0.177118479974329 lpclm = 7.267040315538453E-7
+ wpclm = 6.203018240388111E-7 ppclm = -3.604912502372409E-13 pdiblc1 = 0.242749290147124
+ lpdiblc1 = 2.979647564014913E-7 wpdiblc1 = 4.970203811801911E-7 ppdiblc1 = -1.00573068172574E-12
+ pdiblc2 = -2.185113281247999E-4 lpdiblc2 = 6.637643145622951E-10 wpdiblc2 = 6.363660079716785E-10
+ ppdiblc2 = -6.513333364791723E-16 pdiblcb = -0.025 drout = 0.12432331263201
+ ldrout = 8.816004904228752E-7 wdrout = -1.439733330663757E-8 pdrout = 2.913329189264725E-14
+ pscbe1 = 8.008250796488913E8 lpscbe1 = 6.034187455016056 wpscbe1 = -2.459786855009492
+ ppscbe1 = -1.798955410239063E-5 pscbe2 = -1.16724094431636E-8 lpscbe2 = 2.150883333602323E-14
+ wpscbe2 = 2.080584109298226E-14 ppscbe2 = -2.146131983233702E-20 pvag = 0
+ delta = 0.01 fprout = 0 pdits = 0
+ pditsl = 0 pditsd = 0 lambda = 0
+ vtl = 0 lc = 5E-9 xn = 3
+ alpha0 = 1E-10 alpha1 = 1E-10 beta0 = 7.197826553266499
+ lbeta0 = 2.310234669756333E-6 wbeta0 = -1.310501484340619E-6 pbeta0 = -4.5319440311909E-13
+ aigbacc = 0.43 bigbacc = 0.054 cigbacc = 0.075
+ nigbacc = 1 aigbinv = 0.35 bigbinv = 0.03
+ cigbinv = 6E-3 eigbinv = 1.1 nigbinv = 3
+ aigc = 0.43 bigc = 0.054 cigc = 0.075
+ aigsd = 0.43 bigsd = 0.054 cigsd = 0.075
+ dlcig = 0 nigc = 1 poxedge = 1
+ pigcd = 1 ntox = 1 toxref = 4.23E-9
+ agidl = 2.748348716212996E-10 lagidl = -3.838632912472942E-16 wagidl = -5.212303073881753E-16
+ pagidl = 1.144400882023403E-21 bgidl = 1.401907270501351E9 lbgidl = -47.4690277740255
+ wbgidl = -394.38035113940174 pbgidl = 4.658002782187354E-5 cgidl = 300
+ egidl = 0.1 noia = 1.2E41 noib = 2E25
+ noic = 0 em = 4.1E7 af = 1
+ ef = 0.88 kf = 0 lintnoi = -6E-8
+ tnoia = 1.5 tnoib = 3.5 ntnoi = 1
+ rnoia = 0.577 rnoib = 0.37 xpart = 0
+ cgso = {5.932020000000001E-11/sw_func_tox_lv_ratio} cgdo = {5.932020000000001E-11/sw_func_tox_lv_ratio} cgbo = {0/sw_func_tox_lv_ratio}
+ ckappas = 0.6 cf = 1.2E-11 clc = 1E-7
+ cle = 0.6 dlc = -2.56E-9 dwc = 0
+ vfbcv = -0.1446893 noff = 4 voffcv = -0.1375
+ acde = 0.552 moin = 14.504 cgsl = {7.513892E-12/sw_func_tox_lv_ratio}
+ cgdl = {7.513892E-12/sw_func_tox_lv_ratio} ijthsrev = 0.1 ijthsfwd = 0.1
+ xjbvs = 1 bvs = 12.8 jss = 2.17E-5
+ jsws = 8.200000000000001E-10 cjs = {7.433E-04*sw_func_psd_nw_cj} mjs = 0.34629
+ mjsws = 0.26859 cjsws = {9.2435E-11*sw_func_psd_nw_cj} cjswgs = {2.4701E-10*sw_func_psd_nw_cj}
+ mjswgs = 0.70393 pbs = 0.6587 pbsws = 0.7418
+ pbswgs = 1.3925 xrcrg1 = 12 xrcrg2 = 1
+ rbpb = 50 rbpd = 50 rbps = 50
+ rbdb = 50 rbsb = 50 gbmin = 1E-12
+ tnom = 30 ute = -0.459203677029707 lute = 9.963645903382484E-7
+ wute = 1.369011064625707E-6 pute = -2.97043385496689E-12 kt1 = -0.436825394272762
+ lkt1 = -3.326279003640469E-8 wkt1 = -2.130465293814401E-8 pkt1 = 1.202243190302783E-14
+ kt1l = 0 kt2 = -0.063041029922061 lkt2 = 3.18922223081991E-8
+ wkt2 = 6.659666016480536E-9 pkt2 = -2.356637918979096E-14 ua1 = 1.210171668135681E-9
+ lua1 = 2.645428718002883E-15 wua1 = 4.834100966575749E-15 pua1 = -9.191398802005433E-21
+ ub1 = -1.852125284548357E-19 lub1 = -2.331715943256481E-24 wub1 = -4.009199583771214E-24
+ pub1 = 7.476341669132828E-30 uc1 = 2.973922513190508E-10 luc1 = -4.85015578982596E-16
+ wuc1 = -4.179798748455254E-16 puc1 = 6.72266590081052E-22 at = 4.820118057352592E4
+ lat = 0.076277804098685 wat = 0.047916528427574 pat = -1.102732271093468E-7
+ prt = 0 njs = 1.2556 xtis = 2
+ tpb = 1.9551E-3 tpbsw = 1.4242E-4 tpbswg = 0
+ tcj = 1.2407E-3 tcjsw = 0 tcjswg = 2E-12
+ tvoff = 0 tvfbsdoff = 0 saref = 3E-6
+ sbref = 3E-6 wlod = 0 ku0 = 4.5E-8
+ kvsat = 0.4 kvth0 = 2.65E-8 tku0 = 0
+ llodku0 = 0 wlodku0 = 1 llodvth = 0
+ wlodvth = 1 lku0 = 0 wku0 = 2.5E-7
+ pku0 = 0 lkvth0 = 0 wkvth0 = 2.5E-7
+ pkvth0 = 0 stk2 = 0 lodk2 = 1
+ steta0 = 0 lodeta0 = 1

.model phighvt_model.29 pmos
+ level = 54 lmin = 5E-7 lmax = 1E-6 wmin = 1E-6
+ wmax = 3E-6 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 4.23E-9
+ toxm = 4.23E-9 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 9.999999999999999E22 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {9.364E-9+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {-1.176E-8-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = -5.722E-9 dwb = -1.7864E-8 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = -1.118990379966535 lvth0 = 3.763498445545558E-8
+ wvth0 = 2.548000429398828E-8 pvth0 = -1.543595051501042E-14 k1 = 0.230485385267398
+ lk1 = 1.908927830979374E-7 wk1 = 2.805095778453203E-7 pk1 = -1.874793628780276E-13
+ k2 = 0.085753900930436 lk2 = -5.598229993522777E-8 wk2 = -9.58226110763666E-8
+ pk2 = 6.032246665890886E-14 k3 = -13.778 k3b = 2
+ w0 = 0 lpe0 = 0 lpeb = 0
+ vbm = -3 dvtp0 = 0 dvtp1 = 0
+ dvt0 = 4.05 dvt1 = 0.3 dvt2 = 0.03
+ dvt0w = -4.254 dvt1w = 1.1472E6 dvt2w = -8.96E-3
+ vfbsdoff = 0 u0 = 0.012155474918943 lu0 = -3.560386376854932E-9
+ wu0 = -2.216230325829551E-9 pu0 = 1.840598214235559E-15 ua = -1.320106251996358E-10
+ lua = -6.177488450447711E-16 wua = -4.051508728635674E-16 pua = 2.517876407609994E-22
+ ub = 7.489083458080204E-19 lub = 1.120857073900105E-25 wub = 1.106463108495368E-25
+ pub = 9.4739604104748E-32 uc = -4.767834381684548E-11 luc = 7.652598125261607E-18
+ wuc = -5.269245343295107E-17 puc = 2.929708984413123E-23 ud = 0
+ up = 0 lp = 1 eu = 1.67
+ vsat = 1.210609565054153E5 lvsat = -0.046027506593717 wvsat = -0.124729837830873
+ pvsat = 9.882740659424067E-8 a0 = 1.222347748106977 la0 = 9.727643553470267E-8
+ wa0 = -1.049284098420159E-8 pa0 = -3.498284051577684E-13 ags = -0.163315523851646
+ lags = 7.421620385471018E-7 wags = 1.117664556458961E-7 pags = -6.073268710749804E-14
+ b0 = 0 b1 = 0 keta = 0.021998193129997
+ lketa = -3.84764334290236E-8 wketa = -1.034275525813597E-8 pketa = 1.249335096318091E-14
+ a1 = 0 a2 = 0.384630662716756 la2 = 3.24703672352146E-7
+ wa2 = 6.140267679250918E-7 pa2 = -3.290441717965517E-13 rdsw = 531.92
+ rdswmin = 0 rdw = 0 rdwmin = 0
+ rsw = 0 rswmin = 0 prwb = -0.32348
+ prwg = 0.02 wr = 1 voff = -0.231177336481953
+ lvoff = 2.660728112335513E-8 wvoff = 3.144162127645653E-8 pvoff = -3.077145260722075E-14
+ voffl = 0 minv = 0 nfactor = -0.078623498139761
+ lnfactor = 1.845677923098764E-6 wnfactor = 1.841780880992064E-6 pnfactor = -1.701248130014881E-12
+ eta0 = 0.57950102827249 leta0 = -3.694890233331778E-7 weta0 = -6.301746724326025E-7
+ peta0 = 6.465002103656959E-13 etab = -1.711206322137931 letab = 8.956212452784189E-7
+ wetab = 2.084525710083657E-8 petab = -1.100879056898838E-14 dsub = 0.02217498114864
+ ldsub = 7.013310830494558E-7 wdsub = 1.268807063858322E-6 pdsub = -1.228958801432993E-12
+ cit = 1E-5 cdsc = 0 cdscb = 0
+ cdscd = 0 pclm = -2.485558210621797E-3 lpclm = 5.479637434702553E-7
+ wpclm = 1.593039599296205E-6 ppclm = -1.356107817968688E-12 pdiblc1 = -0.462257479606055
+ lpdiblc1 = 1.019553285379265E-6 wpdiblc1 = 5.206377036319255E-7 ppdiblc1 = -1.02990348360154E-12
+ pdiblc2 = -6.873133926652655E-4 lpdiblc2 = 1.143592603660752E-9 wpdiblc2 = 1.496947288599249E-9
+ ppdiblc2 = -1.532155488827103E-15 pdiblcb = -0.060687498838152 lpdiblcb = 3.652686881082535E-8
+ wpdiblcb = 2.939822022787579E-8 ppdiblcb = -3.008966636763543E-14 drout = 1.015565781195223
+ ldrout = -3.060400100094453E-8 wdrout = -1.52742652449989E-8 pdrout = 3.003084927019884E-14
+ pscbe1 = 8.274072142682632E8 lpscbe1 = -21.173158970603495 wpscbe1 = -54.40862386844437
+ ppscbe1 = 3.518111955760023E-5 pscbe2 = 9.498250122268118E-9 lpscbe2 = -1.597601423874413E-16
+ wpscbe2 = -4.710208779221184E-16 ppscbe2 = 3.159739321230234E-22 pvag = 0
+ delta = 0.01 fprout = 0 pdits = 0
+ pditsl = 0 pditsd = 0 lambda = 0
+ vtl = 0 lc = 5E-9 xn = 3
+ alpha0 = 1E-10 alpha1 = 1E-10 beta0 = 9.363826061282273
+ lbeta0 = 9.329085331202916E-8 wbeta0 = -2.776903385903532E-6 pbeta0 = 1.047697271168583E-12
+ aigbacc = 0.43 bigbacc = 0.054 cigbacc = 0.075
+ nigbacc = 1 aigbinv = 0.35 bigbinv = 0.03
+ cigbinv = 6E-3 eigbinv = 1.1 nigbinv = 3
+ aigc = 0.43 bigc = 0.054 cigc = 0.075
+ aigsd = 0.43 bigsd = 0.054 cigsd = 0.075
+ dlcig = 0 nigc = 1 poxedge = 1
+ pigcd = 1 ntox = 1 toxref = 4.23E-9
+ agidl = -2.622780230873645E-10 lagidl = 1.658824987449176E-16 wagidl = 1.080049326445713E-15
+ pagidl = -4.94540848798258E-22 bgidl = 1.422419293943037E9 lbgidl = -68.46349400705938
+ wbgidl = -414.5082254060713 pbgidl = 6.718130969129517E-5 cgidl = 300
+ egidl = 0.1 noia = 1.2E41 noib = 2E25
+ noic = 0 em = 4.1E7 af = 1
+ ef = 0.88 kf = 0 lintnoi = -6E-8
+ tnoia = 1.5 tnoib = 3.5 ntnoi = 1
+ rnoia = 0.577 rnoib = 0.37 xpart = 0
+ cgso = {5.932020000000001E-11/sw_func_tox_lv_ratio} cgdo = {5.932020000000001E-11/sw_func_tox_lv_ratio} cgbo = {0/sw_func_tox_lv_ratio}
+ ckappas = 0.6 cf = 1.2E-11 clc = 1E-7
+ cle = 0.6 dlc = -2.56E-9 dwc = 0
+ vfbcv = -0.1446893 noff = 4 voffcv = -0.1375
+ acde = 0.552 moin = 14.504 cgsl = {7.513892E-12/sw_func_tox_lv_ratio}
+ cgdl = {7.513892E-12/sw_func_tox_lv_ratio} ijthsrev = 0.1 ijthsfwd = 0.1
+ xjbvs = 1 bvs = 12.8 jss = 2.17E-5
+ jsws = 8.200000000000001E-10 cjs = {7.433E-04*sw_func_psd_nw_cj} mjs = 0.34629
+ mjsws = 0.26859 cjsws = {9.2435E-11*sw_func_psd_nw_cj} cjswgs = {2.4701E-10*sw_func_psd_nw_cj}
+ mjswgs = 0.70393 pbs = 0.6587 pbsws = 0.7418
+ pbswgs = 1.3925 xrcrg1 = 12 xrcrg2 = 1
+ rbpb = 50 rbpd = 50 rbps = 50
+ rbdb = 50 rbsb = 50 gbmin = 1E-12
+ tnom = 30 ute = 0.981937780010695 lute = -4.786725137717428E-7
+ wute = -2.864993388590444E-6 pute = 1.363154382988904E-12 kt1 = -0.4701530672535
+ lkt1 = 8.487498128403E-10 wkt1 = 5.187906040586006E-8 pkt1 = -6.28825623788272E-14
+ kt1l = 0 kt2 = -7.750059266772795E-3 lkt2 = -2.469919197690102E-8
+ wkt2 = -5.637502333480736E-8 pkt2 = 4.095088605503922E-14 ua1 = 5.728924778387321E-9
+ lua1 = -1.979605465401874E-15 wua1 = -9.123089027094664E-15 pua1 = 5.094064300316106E-21
+ ub1 = -3.683235567602748E-18 lub1 = 1.24858059777219E-24 wub1 = 7.917308573706308E-24
+ pub1 = -4.730677960208565E-30 uc1 = -3.519863943457512E-10 luc1 = 1.796364524282422E-16
+ wuc1 = 6.805024576894275E-16 puc1 = -4.520520469151228E-22 at = 2.146257009906882E5
+ lat = -0.094061021038689 wat = -0.12259877270393 pat = 6.42525939047704E-8
+ prt = 0 njs = 1.2556 xtis = 2
+ tpb = 1.9551E-3 tpbsw = 1.4242E-4 tpbswg = 0
+ tcj = 1.2407E-3 tcjsw = 0 tcjswg = 2E-12
+ tvoff = 0 tvfbsdoff = 0 saref = 2.75E-6
+ sbref = 2.74E-6 wlod = 0 ku0 = 4.5E-8
+ kvsat = 0.4 kvth0 = 2.65E-8 tku0 = 0
+ llodku0 = 0 wlodku0 = 1 llodvth = 0
+ wlodvth = 1 lku0 = 0 wku0 = 2.5E-7
+ pku0 = 0 lkvth0 = 0 wkvth0 = 2.5E-7
+ pkvth0 = 0 stk2 = 0 lodk2 = 1
+ steta0 = 0 lodeta0 = 1

.model phighvt_model.30 pmos
+ level = 54 lmin = 2.5E-7 lmax = 5E-7 wmin = 1E-6
+ wmax = 3E-6 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 4.23E-9
+ toxm = 4.23E-9 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 9.999999999999999E22 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {9.364E-9+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {-1.176E-8-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = -5.722E-9 dwb = -1.7864E-8 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = -1.036351339792998 lvth0 = -5.62820585619407E-9
+ wvth0 = -1.687463560121697E-8 pvth0 = 6.737550562927434E-15 k1 = 0.432704164917531
+ lk1 = 8.502720757549985E-8 wk1 = 5.995203713860133E-8 pk1 = -7.201307916724604E-14
+ k2 = 0.031233527024181 lk2 = -2.743979378782474E-8 wk2 = -3.17066854501418E-8
+ pk2 = 2.675649727506765E-14 k3 = -13.778 k3b = 2
+ w0 = 0 lpe0 = 0 lpeb = 0
+ vbm = -3 dvtp0 = 0 dvtp1 = 0
+ dvt0 = 4.05 dvt1 = 0.3 dvt2 = 0.03
+ dvt0w = -4.254 dvt1w = 1.1472E6 dvt2w = -8.96E-3
+ vfbsdoff = 0 u0 = 5.414750141161794E-3 lu0 = -3.148214119098022E-11
+ wu0 = 1.970281421997059E-9 pu0 = -3.511244159866286E-16 ua = -9.47278183247948E-10
+ lua = -1.909399730553187E-16 wua = -2.787066885207248E-16 pua = 1.855915813738345E-22
+ ub = 3.939603561701322E-19 lub = 2.979080789252377E-25 wub = 8.555311242321744E-25
+ pub = -2.952224933973304E-31 uc = -3.735917830284466E-11 luc = 2.250308595371896E-18
+ wuc = -2.448077287861522E-17 puc = 1.452771084032533E-23 ud = 0
+ up = 0 lp = 1 eu = 1.67
+ vsat = -1.023326618887403E4 lvsat = 0.022707644871198 wvsat = 0.107268837951654
+ pvsat = -2.262854015142805E-8 a0 = 2.001776910118605 la0 = -3.107703193616248E-7
+ wa0 = -1.128745778158217E-6 pa0 = 2.355993725115723E-13 ags = -0.242868114125184
+ lags = 7.838094106071045E-7 wags = 1.166881076718472E-6 pags = -6.131062935314129E-13
+ b0 = 0 b1 = 0 keta = -0.016001093926732
+ lketa = -1.85830466690852E-8 wketa = -2.604042970369088E-8 pketa = 2.071139748891782E-14
+ a1 = 0 a2 = 1.228998067590488 la2 = -1.173395514473504E-7
+ wa2 = -3.035551300963066E-8 pa2 = 8.302839918394176E-15 rdsw = 531.92
+ rdswmin = 0 rdw = 0 rdwmin = 0
+ rsw = 0 rswmin = 0 prwb = -0.32348
+ prwg = 0.02 wr = 1 voff = -0.116215518800203
+ lvoff = -3.357752966939426E-8 wvoff = -8.102257717273758E-8 pvoff = 2.810580456490135E-14
+ voffl = 0 minv = 0 nfactor = 5.64599978316097
+ lnfactor = -1.151276857127794E-6 wnfactor = -4.017800962902757E-6 pnfactor = 1.366360156900936E-12
+ eta0 = -0.800533780047856 leta0 = 3.529867995186895E-7 weta0 = 1.26636466341512E-6
+ peta0 = -3.463760627373034E-13 etab = 9.798797891017309E-5 letab = -2.807871539495105E-10
+ wetab = -1.373731715705143E-9 petab = 6.232944562475613E-16 dsub = 2.332982177378136
+ ldsub = -5.084227003206105E-7 wdsub = -2.623756309091292E-6 pdsub = 8.088759755735886E-13
+ cit = 1E-5 cdsc = 0 cdscb = 0
+ cdscd = 0 pclm = 1.487984056056094 lpclm = -2.323269089906557E-7
+ wpclm = -2.088472986552131E-6 ppclm = 5.712376509746321E-13 pdiblc1 = 2.714325191814697
+ lpdiblc1 = -6.434512747629265E-7 wpdiblc1 = -3.079765725866971E-6 ppdiblc1 = 8.549797198097227E-13
+ pdiblc2 = -5.003693753443018E-3 lpdiblc2 = 3.403304050135121E-9 wpdiblc2 = -4.877494151530442E-9
+ ppdiblc2 = 1.804992093909592E-15 pdiblcb = -0.056414444942174 lpdiblcb = 3.428983963520278E-8
+ wpdiblcb = 2.476468467183228E-7 ppdiblcb = -1.443471873079142E-13 drout = 1.551807682972029
+ ldrout = -3.113373614191379E-7 wdrout = 7.060755340660586E-9 pdrout = 1.833801929319439E-14
+ pscbe1 = 7.729250162838502E8 lpscbe1 = 7.349361318196452 wpscbe1 = 26.599003853633366
+ ppscbe1 = -7.227993707461904E-6 pscbe2 = 9.257822908086217E-9 lpscbe2 = -3.389168721893256E-17
+ wpscbe2 = 2.550236571112633E-16 ppscbe2 = -6.412490285765253E-23 pvag = 0
+ delta = 0.01 fprout = 0 pdits = 0
+ pditsl = 0 pditsd = 0 lambda = 0
+ vtl = 0 lc = 5E-9 xn = 3
+ alpha0 = 1E-10 alpha1 = 1E-10 beta0 = 10.573525466633852
+ lbeta0 = -5.400109793776305E-7 wbeta0 = -2.008029813310324E-6 pbeta0 = 6.451765784445864E-13
+ aigbacc = 0.43 bigbacc = 0.054 cigbacc = 0.075
+ nigbacc = 1 aigbinv = 0.35 bigbinv = 0.03
+ cigbinv = 6E-3 eigbinv = 1.1 nigbinv = 3
+ aigc = 0.43 bigc = 0.054 cigc = 0.075
+ aigsd = 0.43 bigsd = 0.054 cigsd = 0.075
+ dlcig = 0 nigc = 1 poxedge = 1
+ pigcd = 1 ntox = 1 toxref = 4.23E-9
+ agidl = 4.8908323928826E-12 lagidl = 2.601425952389875E-17 wagidl = 2.835462983304061E-16
+ pagidl = -7.755558351933267E-23 bgidl = 1.685496056929084E9 lbgidl = -206.18944096551493
+ wbgidl = -952.1864786991808 pbgidl = 3.486666288553038E-4 cgidl = 300
+ egidl = 0.1 noia = 1.2E41 noib = 2E25
+ noic = 0 em = 4.1E7 af = 1
+ ef = 0.88 kf = 0 lintnoi = -6E-8
+ tnoia = 1.5 tnoib = 3.5 ntnoi = 1
+ rnoia = 0.577 rnoib = 0.37 xpart = 0
+ cgso = {5.932020000000001E-11/sw_func_tox_lv_ratio} cgdo = {5.932020000000001E-11/sw_func_tox_lv_ratio} cgbo = {0/sw_func_tox_lv_ratio}
+ ckappas = 0.6 cf = 1.2E-11 clc = 1E-7
+ cle = 0.6 dlc = -2.56E-9 dwc = 0
+ vfbcv = -0.1446893 noff = 4 voffcv = -0.1375
+ acde = 0.552 moin = 14.504 cgsl = {7.513892E-12/sw_func_tox_lv_ratio}
+ cgdl = {7.513892E-12/sw_func_tox_lv_ratio} ijthsrev = 0.1 ijthsfwd = 0.1
+ xjbvs = 1 bvs = 12.8 jss = 2.17E-5
+ jsws = 8.200000000000001E-10 cjs = {7.433E-04*sw_func_psd_nw_cj} mjs = 0.34629
+ mjsws = 0.26859 cjsws = {9.2435E-11*sw_func_psd_nw_cj} cjswgs = {2.4701E-10*sw_func_psd_nw_cj}
+ mjswgs = 0.70393 pbs = 0.6587 pbsws = 0.7418
+ pbswgs = 1.3925 xrcrg1 = 12 xrcrg2 = 1
+ rbpb = 50 rbpd = 50 rbps = 50
+ rbdb = 50 rbsb = 50 gbmin = 1E-12
+ tnom = 30 ute = -0.322288835129263 lute = 2.041162037863281E-7
+ wute = 8.359702386882896E-7 pute = -5.743740951640585E-13 kt1 = -0.461482314362547
+ lkt1 = -3.690562740631326E-9 wkt1 = -9.733836021117772E-8 pkt1 = 1.523574166260437E-14
+ kt1l = 0 kt2 = -0.062079437560823 lkt2 = 3.743324147600199E-9
+ wkt2 = 5.067738325226774E-8 pkt2 = -1.509318984142633E-14 ua1 = 1.330866595791479E-9
+ lua1 = 3.228659543507009E-16 wua1 = 3.656071484238083E-15 pua1 = -1.596081810576813E-21
+ ub1 = -4.571458113931081E-19 lub1 = -4.403419113986803E-25 wub1 = -4.375616599821293E-24
+ pub1 = 1.704914226636604E-30 uc1 = 1.172374923074039E-10 luc1 = -6.601163671241754E-17
+ wuc1 = -4.051396285068132E-16 puc1 = 1.16303298050333E-22 at = 4.032802764631296E4
+ lat = -2.81270308944128E-3 wat = -0.044825667750906 pat = 2.35368179997634E-8
+ prt = 0 njs = 1.2556 xtis = 2
+ tpb = 1.9551E-3 tpbsw = 1.4242E-4 tpbswg = 0
+ tcj = 1.2407E-3 tcjsw = 0 tcjswg = 2E-12
+ tvoff = 0 tvfbsdoff = 0 saref = 1.75E-6
+ sbref = 1.74E-6 wlod = 0 ku0 = 4.5E-8
+ kvsat = 0.4 kvth0 = 2.65E-8 tku0 = 0
+ llodku0 = 0 wlodku0 = 1 llodvth = 0
+ wlodvth = 1 lku0 = 0 wku0 = 2.5E-7
+ pku0 = 0 lkvth0 = 0 wkvth0 = 2.5E-7
+ pkvth0 = 0 stk2 = 0 lodk2 = 1
+ steta0 = 0 lodeta0 = 1

.model phighvt_model.31 pmos
+ level = 54 lmin = 1.8E-7 lmax = 2.5E-7 wmin = 1E-6
+ wmax = 3E-6 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 4.23E-9
+ toxm = 4.23E-9 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 9.999999999999999E22 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {9.364E-9+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {-1.176E-8-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = -5.722E-9 dwb = -1.7864E-8 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = -0.978491680691551 lvth0 = -2.1453979813622E-8
+ wvth0 = -3.986122366453228E-8 pvth0 = 1.302484213000544E-14 k1 = 0.085401790352232
+ lk1 = 1.800213530666004E-7 wk1 = -7.20715530328475E-7 pk1 = 1.415151138863486E-13
+ k2 = 0.223483693247248 lk2 = -8.002405925315811E-8 wk2 = 1.915114723177419E-7
+ pk2 = -3.429813323760389E-14 k3 = -13.778 k3b = 2
+ w0 = 0 lpe0 = 0 lpeb = 0
+ vbm = -3 dvtp0 = 0 dvtp1 = 0
+ dvt0 = 4.05 dvt1 = 0.3 dvt2 = 0.03
+ dvt0w = -4.254 dvt1w = 1.1472E6 dvt2w = -8.96E-3
+ vfbsdoff = 0 u0 = 7.989256064291428E-3 lu0 = -7.356610012853982E-10
+ wu0 = 8.171400260508971E-9 pu0 = -2.047254440696406E-15 ua = -8.518349483012087E-10
+ lua = -2.170456066779507E-16 wua = 3.133476820696168E-15 pua = -7.477088520671701E-22
+ ub = 8.033482526153999E-19 lub = 1.859323014895282E-25 wub = -2.12906697709323E-24
+ pub = 5.21124779277194E-31 uc = -9.177597757938408E-11 luc = 1.713439153349096E-17
+ wuc = 1.182855337344049E-16 puc = -2.452172934446792E-23 ud = 0
+ up = 0 lp = 1 eu = 1.67
+ vsat = -2.37557222092626E3 lvsat = 0.020558408417085 wvsat = -0.075165225944239
+ pvsat = 2.72708250053766E-8 a0 = 1.40276047357184 la0 = -1.469273436373538E-7
+ wa0 = -1.714554107788868E-6 pa0 = 3.958296668321478E-13 ags = 6.614001771879774
+ lags = -1.091681640612972E-6 wags = -4.199156877533952E-6 pags = 8.5461240771571E-13
+ b0 = 0 b1 = 0 keta = -0.084000741279438
+ lketa = 1.621687482699754E-11 wketa = 9.991477100043185E-8 pketa = -1.373986900767383E-14
+ a1 = 0 a2 = 1.065523986242529 la2 = -7.262612071705655E-8
+ wa2 = 3.969817764973988E-7 pa2 = -1.085824555075685E-13 rdsw = 531.92
+ rdswmin = 0 rdw = 0 rdwmin = 0
+ rsw = 0 rswmin = 0 prwb = -0.32348
+ prwg = 0.02 wr = 1 voff = -0.201576546096548
+ lvoff = -1.022958148329822E-8 wvoff = 1.372157394643679E-7 pvoff = -3.158673980167974E-14
+ voffl = 0 minv = 0 nfactor = -0.475222239757528
+ lnfactor = 5.229997905808733E-7 wnfactor = 4.752053767601366E-6 pnfactor = -1.032370508986552E-12
+ eta0 = 0.372620728994316 leta0 = 3.210557820547457E-8 weta0 = 3.499395340296564E-7
+ peta0 = -9.57154613477916E-14 etab = -9.285810249999998E-4 wetab = 9.050576095637997E-10
+ dsub = 0.842292208820679 ldsub = -1.006891801207745E-7 wdsub = -5.581843728768861E-7
+ pdsub = 2.439007395802242E-13 cit = 1E-5 cdsc = 0
+ cdscb = 0 cdscd = 0 pclm = 0.286343155740852
+ lpclm = 9.634591006356946E-8 wpclm = 2.171123389471958E-7 ppclm = -5.938604725594365E-14
+ pdiblc1 = -0.018226450790969 lpdiblc1 = 1.039562505225749E-7 wpdiblc1 = 4.489805093777009E-7
+ ppdiblc1 = -1.102029504543998E-13 pdiblc2 = 4.272437443945823E-4 lpdiblc2 = 1.91783402572658E-9
+ wpdiblc2 = 6.477059951619321E-9 ppdiblc2 = -1.30070554438393E-15 pdiblcb = 1.052243915311513
+ lpdiblcb = -2.689503950613855E-7 wpdiblcb = -1.481315805250139E-6 ppdiblcb = 3.285586772584994E-13
+ drout = -0.651928392658716 ldrout = 2.914285299873836E-7 wdrout = 1.118193982415284E-6
+ pdrout = -2.855791409762566E-13 pscbe1 = 7.9997105E8 pscbe2 = 4.793980044031212E-9
+ lpscbe2 = 1.187058612957392E-15 wpscbe2 = 1.140613084791645E-14 ppscbe2 = -3.114175741686685E-21
+ pvag = 0 delta = 0.01 fprout = 0
+ pdits = 0 pditsl = 0 pditsd = 0
+ lambda = 0 vtl = 0 lc = 5E-9
+ xn = 3 alpha0 = 1E-10 alpha1 = 1E-10
+ beta0 = 8.031909947876862 lbeta0 = 1.551716973127818E-7 wbeta0 = 5.267241866010946E-8
+ pbeta0 = 8.153330395603338E-14 aigbacc = 0.43 bigbacc = 0.054
+ cigbacc = 0.075 nigbacc = 1 aigbinv = 0.35
+ bigbinv = 0.03 cigbinv = 6E-3 eigbinv = 1.1
+ nigbinv = 3 aigc = 0.43 bigc = 0.054
+ cigc = 0.075 aigsd = 0.43 bigsd = 0.054
+ cigsd = 0.075 dlcig = 0 nigc = 1
+ poxedge = 1 pigcd = 1 ntox = 1
+ toxref = 4.23E-9 agidl = -6.780057631718106E-10 lagidl = 2.128001363427536E-16
+ wagidl = 4.077555285204408E-16 pagidl = -1.115292921609109E-22 bgidl = 7.329634360818298E8
+ lbgidl = 54.347281488625946 wbgidl = 1.260351188592914E3 pbgidl = -2.565066739024298E-4
+ cgidl = 300 egidl = 0.1 noia = 1.2E41
+ noib = 2E25 noic = 0 em = 4.1E7
+ af = 1 ef = 0.88 kf = 0
+ lintnoi = -6E-8 tnoia = 1.5 tnoib = 3.5
+ ntnoi = 1 rnoia = 0.577 rnoib = 0.37
+ xpart = 0 cgso = {5.932020000000001E-11/sw_func_tox_lv_ratio} cgdo = {5.932020000000001E-11/sw_func_tox_lv_ratio}
+ cgbo = {0/sw_func_tox_lv_ratio} ckappas = 0.6 cf = 1.2E-11
+ clc = 1E-7 cle = 0.6 dlc = -2.56E-9
+ dwc = 0 vfbcv = -0.1446893 noff = 4
+ voffcv = -0.1375 acde = 0.552 moin = 14.504
+ cgsl = {7.513892E-12/sw_func_tox_lv_ratio} cgdl = {7.513892E-12/sw_func_tox_lv_ratio} ijthsrev = 0.1
+ ijthsfwd = 0.1 xjbvs = 1 bvs = 12.8
+ jss = 2.17E-5 jsws = 8.200000000000001E-10 cjs = {7.433E-04*sw_func_psd_nw_cj}
+ mjs = 0.34629 mjsws = 0.26859 cjsws = {9.2435E-11*sw_func_psd_nw_cj}
+ cjswgs = {2.4701E-10*sw_func_psd_nw_cj} mjswgs = 0.70393 pbs = 0.6587
+ pbsws = 0.7418 pbswgs = 1.3925 xrcrg1 = 12
+ xrcrg2 = 1 rbpb = 50 rbpd = 50
+ rbps = 50 rbdb = 50 rbsb = 50
+ gbmin = 1E-12 tnom = 30 ute = 1.389962163503255
+ lute = -2.642186893596385E-7 wute = -3.970498571271679E-6 pute = 7.402912537361917E-13
+ kt1 = -0.388143259089646 lkt1 = -2.375026113887521E-8 wkt1 = -6.700231554098271E-8
+ pkt1 = 6.938226724412629E-15 kt1l = 0 kt2 = -0.038980561350907
+ lkt2 = -2.57468047333602E-9 wkt2 = -4.22094188076631E-8 pkt2 = 1.031320825800595E-14
+ ua1 = 6.391767302714457E-9 lua1 = -1.061391607006872E-15 wua1 = -5.713745054536837E-15
+ pua1 = 9.66750409108903E-22 ub1 = -5.518115788225166E-18 lub1 = 9.439345966644243E-25
+ wub1 = 3.696700749545094E-24 pub1 = -5.030260147620897E-31 uc1 = -4.212586141027812E-10
+ luc1 = 8.127781831289626E-17 wuc1 = 1.162369981311315E-16 puc1 = -2.63036368676776E-23
+ at = 1.476361858519754E5 lat = -0.032163630521854 wat = -0.014617841822889
+ pat = 1.527437345193208E-8 prt = 0 njs = 1.2556
+ xtis = 2 tpb = 1.9551E-3 tpbsw = 1.4242E-4
+ tpbswg = 0 tcj = 1.2407E-3 tcjsw = 0
+ tcjswg = 2E-12 tvoff = 0 tvfbsdoff = 0
+ saref = 1.25E-6 sbref = 1.24E-6 wlod = 0
+ ku0 = 4.5E-8 kvsat = 0.4 kvth0 = 2.65E-8
+ tku0 = 0 llodku0 = 0 wlodku0 = 1
+ llodvth = 0 wlodvth = 1 lku0 = 0
+ wku0 = 2.5E-7 pku0 = 0 lkvth0 = 0
+ wkvth0 = 2.5E-7 pkvth0 = 0 stk2 = 0
+ lodk2 = 1 steta0 = 0 lodeta0 = 1

.model phighvt_model.32 pmos
+ level = 54 lmin = 1.5E-7 lmax = 1.8E-7 wmin = 1E-6
+ wmax = 3E-6 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 4.23E-9
+ toxm = 4.23E-9 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 9.999999999999999E22 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {9.364E-9+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {-1.176E-8-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = -5.722E-9 dwb = -1.7864E-8 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = -0.96050049426552 lvth0 = -2.511554607504769E-8
+ wvth0 = 1.637428629933272E-7 pvth0 = -2.841266158660214E-14 k1 = 1.65416942839622
+ lk1 = -1.392542366281121E-7 wk1 = -1.72163694870086E-7 pk1 = 2.987384433385732E-14
+ k2 = -0.630983069317919 lk2 = 9.387701626410459E-8 wk2 = 2.32090269940094E-7
+ pk2 = -4.255673012970498E-14 k3 = -13.778 k3b = 2
+ w0 = 0 lpe0 = 0 lpeb = 0
+ vbm = -3 dvtp0 = 0 dvtp1 = 0
+ dvt0 = 4.05 dvt1 = 0.3 dvt2 = 0.03
+ dvt0w = -4.254 dvt1w = 1.1472E6 dvt2w = -8.96E-3
+ vfbsdoff = 0 u0 = 0.017596375592773 lu0 = -2.690901967721987E-9
+ wu0 = -1.238401688107484E-8 pu0 = 2.136184055958732E-15 ua = 2.311775426792899E-9
+ lua = -8.609035902171038E-16 wua = -3.666121650636188E-15 pua = 6.361454288183913E-22
+ ub = -1.616231746096733E-18 lub = 6.783652228274215E-25 wub = 2.588821696132905E-24
+ pub = -4.390599234977889E-31 uc = -1.050103565928429E-10 luc = 1.98278523503101E-17
+ wuc = -1.494191729472796E-17 puc = 2.592721488981195E-24 ud = 0
+ up = 0 lp = 1 eu = 1.67
+ vsat = 2.108228866227198E5 lvsat = -0.022831741926774 wvsat = 0.399106607373502
+ pvsat = -6.925297851144999E-8 a0 = -2.127217028533755 la0 = 5.71493677591177E-7
+ wa0 = 1.562787160498577E-6 pa0 = -2.711748280897131E-13 ags = 1.25
+ b0 = 0 b1 = 0 keta = -0.338035086632913
+ lketa = 5.171728684116624E-8 wketa = 1.689637399293255E-8 pketa = 3.156035151292429E-15
+ a1 = 0 a2 = 2.190407457300764 la2 = -3.015624047468284E-7
+ wa2 = -9.262908118272619E-7 pa2 = 1.607299816682664E-13 rdsw = 531.92
+ rdswmin = 0 rdw = 0 rdwmin = 0
+ rsw = 0 rswmin = 0 prwb = -0.32348
+ prwg = 0.02 wr = 1 voff = -0.197596599682253
+ lvoff = -1.103958017753552E-8 wvoff = -1.220197501963858E-7 pvoff = 2.117286705407686E-14
+ voffl = 0 minv = 0 nfactor = 3.089329324580707
+ lnfactor = -2.024577437932443E-7 wnfactor = -2.174417540144057E-6 pnfactor = 3.773049315657967E-13
+ eta0 = 0.763884965679928 leta0 = -4.752451924478106E-8 weta0 = -8.165255794025297E-7
+ peta0 = 1.41683518537927E-13 etab = -6.26334367359999E-3 letab = 1.08573089424307E-9
+ wetab = 6.139910823280809E-9 petab = -1.065397326055686E-15 dsub = -1.471988490346329
+ ldsub = 3.70313227773695E-7 wdsub = 4.343301867077337E-6 pdsub = -7.536497399752595E-13
+ cit = 1E-5 cdsc = 0 cdscb = 0
+ cdscd = 0 pclm = 0.372684797118254 lpclm = 7.877365921044046E-8
+ wpclm = -5.066448011136777E-7 ppclm = 8.791300588924535E-14 pdiblc1 = 2.255509707386559
+ lpdiblc1 = -3.587945323897157E-7 wpdiblc1 = -6.275479061950028E-7 ppdiblc1 = 1.088921126829569E-13
+ pdiblc2 = -0.151763080409141 lpdiblc2 = 3.289160879745416E-8 wpdiblc2 = 2.890210573750048E-8
+ ppdiblc2 = -5.864650862726465E-15 pdiblcb = -0.525190447239546 lpdiblcb = 5.208904640500607E-8
+ wpdiblcb = 9.027094857997019E-7 ppdiblcb = -1.566381499759642E-13 drout = -0.481433154083946
+ ldrout = 2.567293390326464E-7 wdrout = -1.933476722503264E-6 pdrout = 3.354968808887662E-13
+ pscbe1 = 8E8 pscbe2 = 1.81986634274208E-8 lpscbe2 = -1.541062549230057E-15
+ wpscbe2 = -2.642666638395763E-14 ppscbe2 = 4.585555150944328E-21 pvag = 0
+ delta = 0.01 fprout = 0 pdits = 0
+ pditsl = 0 pditsd = 0 lambda = 0
+ vtl = 0 lc = 5E-9 xn = 3
+ alpha0 = 1E-10 alpha1 = 1E-10 beta0 = 7.111986328822698
+ lbeta0 = 3.423945522626854E-7 wbeta0 = 3.075106486724623E-6 pbeta0 = -5.335924775764565E-13
+ aigbacc = 0.43 bigbacc = 0.054 cigbacc = 0.075
+ nigbacc = 1 aigbinv = 0.35 bigbinv = 0.03
+ cigbinv = 6E-3 eigbinv = 1.1 nigbinv = 3
+ aigc = 0.43 bigc = 0.054 cigc = 0.075
+ aigsd = 0.43 bigsd = 0.054 cigsd = 0.075
+ dlcig = 0 nigc = 1 poxedge = 1
+ pigcd = 1 ntox = 1 toxref = 4.23E-9
+ agidl = 3.449353077208712E-9 lagidl = -6.271999348514907E-16 wagidl = -7.702144238129276E-15
+ pagidl = 1.53899750834764E-21 bgidl = 1E9 cgidl = 300
+ egidl = 0.1 noia = 1.2E41 noib = 2E25
+ noic = 0 em = 4.1E7 af = 1
+ ef = 0.88 kf = 0 lintnoi = -6E-8
+ tnoia = 1.5 tnoib = 3.5 ntnoi = 1
+ rnoia = 0.577 rnoib = 0.37 xpart = 0
+ cgso = {5.932020000000001E-11/sw_func_tox_lv_ratio} cgdo = {5.932020000000001E-11/sw_func_tox_lv_ratio} cgbo = {0/sw_func_tox_lv_ratio}
+ ckappas = 0.6 cf = 1.2E-11 clc = 1E-7
+ cle = 0.6 dlc = -2.56E-9 dwc = 0
+ vfbcv = -0.1446893 noff = 4 voffcv = -0.1375
+ acde = 0.552 moin = 14.504 cgsl = {7.513892E-12/sw_func_tox_lv_ratio}
+ cgdl = {7.513892E-12/sw_func_tox_lv_ratio} ijthsrev = 0.1 ijthsfwd = 0.1
+ xjbvs = 1 bvs = 12.8 jss = 2.17E-5
+ jsws = 8.200000000000001E-10 cjs = {7.433E-04*sw_func_psd_nw_cj} mjs = 0.34629
+ mjsws = 0.26859 cjsws = {9.2435E-11*sw_func_psd_nw_cj} cjswgs = {2.4701E-10*sw_func_psd_nw_cj}
+ mjswgs = 0.70393 pbs = 0.6587 pbsws = 0.7418
+ pbswgs = 1.3925 xrcrg1 = 12 xrcrg2 = 1
+ rbpb = 50 rbpd = 50 rbps = 50
+ rbdb = 50 rbsb = 50 gbmin = 1E-12
+ tnom = 30 ute = 1.694788743905437 lute = -3.262569950030905E-7
+ wute = -2.999642550081734E-6 pute = 5.427026363036142E-13 kt1 = -0.119314705920001
+ lkt1 = -7.84622482799614E-8 wkt1 = 1.151452687270506E-7 pkt1 = -3.013244962581749E-14
+ kt1l = 0 kt2 = -0.179196542873088 lkt2 = 2.596207608605816E-8
+ wkt2 = 2.773945009955042E-7 pkt2 = -5.473258150033467E-14 ua1 = 6.285408428052469E-9
+ lua1 = -1.039745448835664E-15 wua1 = -6.537032813014461E-15 pua1 = 1.134305933714269E-21
+ ub1 = -6.286066967838709E-18 lub1 = 1.100228020739372E-24 wub1 = 8.31088405951091E-24
+ pub1 = -1.442104602006333E-30 uc1 = 1.888518123566076E-10 luc1 = -4.289185568011854E-17
+ wuc1 = -8.823610026765732E-17 puc1 = 1.531072811844389E-23 at = -4.244454350671254E5
+ lat = 0.084266420967601 wat = 0.515906390743732 pat = -9.269791836002666E-8
+ prt = 0 njs = 1.2556 xtis = 2
+ tpb = 1.9551E-3 tpbsw = 1.4242E-4 tpbswg = 0
+ tcj = 1.2407E-3 tcjsw = 0 tcjswg = 2E-12
+ tvoff = 0 tvfbsdoff = 0 saref = 1.1E-6
+ sbref = 1.1E-6 wlod = 0 ku0 = 4.5E-8
+ kvsat = 0.4 kvth0 = 2.65E-8 tku0 = 0
+ llodku0 = 0 wlodku0 = 1 llodvth = 0
+ wlodvth = 1 lku0 = 0 wku0 = 2.5E-7
+ pku0 = 0 lkvth0 = 0 wkvth0 = 2.5E-7
+ pkvth0 = 0 stk2 = 0 lodk2 = 1
+ steta0 = 0 lodeta0 = 1

.model phighvt_model.33 pmos
+ level = 54 lmin = 8E-6 lmax = 2.02E-5 wmin = 5.5E-7
+ wmax = 1E-6 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 4.23E-9
+ toxm = 4.23E-9 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 9.999999999999999E22 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {9.364E-9+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {-1.176E-8-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = -5.722E-9 dwb = -1.7864E-8 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = -1.100899108531555 wvth0 = 1.24782556325765E-8
+ k1 = 0.440441229602311 wk1 = 6.943932447360951E-9 k2 = 0.016141931735413
+ wk2 = 4.752475222047489E-9 k3 = -13.778 k3b = 2
+ w0 = 0 lpe0 = 0 lpeb = 0
+ vbm = -3 dvtp0 = 0 dvtp1 = 0
+ dvt0 = 4.05 dvt1 = 0.3 dvt2 = 0.03
+ dvt0w = -4.254 dvt1w = 1.1472E6 dvt2w = -8.96E-3
+ vfbsdoff = 0 u0 = 0.01007186173648 wu0 = -1.033438123479201E-9
+ ua = -9.917710680666667E-10 wua = 2.600920587730342E-16 ub = 1.713539570411022E-18
+ wub = -7.146294486844446E-25 uc = -2.998833915823998E-11 wuc = -4.100595350576353E-17
+ ud = 0 up = 0 lp = 1
+ eu = 1.67 vsat = 2.774802639709156E5 wvsat = -0.114975899267268
+ a0 = 1.296014829434667 wa0 = -3.989540833301424E-8 ags = 0.395313352528533
+ wags = -1.49397045382379E-7 b0 = -2.652936247111112E-8 wb0 = 2.603252057075215E-14
+ b1 = -3.447837219555557E-11 wb1 = 3.38326612410772E-17 keta = -0.012496273158164
+ wketa = 1.042706806005747E-8 a1 = 0 a2 = 0.8
+ rdsw = 531.92 rdswmin = 0 rdw = 0
+ rdwmin = 0 rsw = 0 rswmin = 0
+ prwb = -0.32348 prwg = 0.02 wr = 1
+ voff = -0.22219315336 wvoff = 9.972896325633944E-9 voffl = 0
+ minv = 0 nfactor = 2.200787116933333 wnfactor = -3.78853631718606E-7
+ eta0 = 0.08 etab = -0.07 dsub = 0.56
+ cit = 1E-5 cdsc = 0 cdscb = 0
+ cdscd = 0 pclm = 0.14095898 pdiblc1 = 0.39
+ pdiblc2 = 3.052192647758223E-4 wpdiblc2 = 1.381508829633936E-11 pdiblcb = -0.072618336538133
+ wpdiblcb = -8.095611111071285E-8 drout = 0.56 pscbe1 = 8E8
+ pscbe2 = -2.165432053223114E-9 wpscbe2 = 7.448732574411951E-15 pvag = 0
+ delta = 0.01 fprout = 0 pdits = 0
+ pditsl = 0 pditsd = 0 lambda = 0
+ vtl = 0 lc = 5E-9 xn = 3
+ alpha0 = 1E-10 alpha1 = 1E-10 beta0 = 10.149306399088001
+ wbeta0 = -3.798226309256281E-6 aigbacc = 0.43 bigbacc = 0.054
+ cigbacc = 0.075 nigbacc = 1 aigbinv = 0.35
+ bigbinv = 0.03 cigbinv = 6E-3 eigbinv = 1.1
+ nigbinv = 3 aigc = 0.43 bigc = 0.054
+ cigc = 0.075 aigsd = 0.43 bigsd = 0.054
+ cigsd = 0.075 dlcig = 0 nigc = 1
+ poxedge = 1 pigcd = 1 ntox = 1
+ toxref = 4.23E-9 agidl = 3.369193107429333E-10 wagidl = 1.061524538212203E-16
+ bgidl = 1E9 cgidl = 300 egidl = 1.812754997677333
+ wegidl = -9.099387731260325E-7 noia = 1.2E41 noib = 2E25
+ noic = 0 em = 4.1E7 af = 1
+ ef = 0.88 kf = 0 lintnoi = -6E-8
+ tnoia = 1.5 tnoib = 3.5 ntnoi = 1
+ rnoia = 0.577 rnoib = 0.37 xpart = 0
+ cgso = {5.932020000000001E-11/sw_func_tox_lv_ratio} cgdo = {5.932020000000001E-11/sw_func_tox_lv_ratio} cgbo = {0/sw_func_tox_lv_ratio}
+ ckappas = 0.6 cf = 1.2E-11 clc = 1E-7
+ cle = 0.6 dlc = -2.56E-9 dwc = 0
+ vfbcv = -0.1446893 noff = 4 voffcv = -0.1375
+ acde = 0.552 moin = 14.504 cgsl = {7.513892E-12/sw_func_tox_lv_ratio}
+ cgdl = {7.513892E-12/sw_func_tox_lv_ratio} ijthsrev = 0.1 ijthsfwd = 0.1
+ xjbvs = 1 bvs = 12.8 jss = 2.17E-5
+ jsws = 8.200000000000001E-10 cjs = {7.433E-04*sw_func_psd_nw_cj} mjs = 0.34629
+ mjsws = 0.26859 cjsws = {9.2435E-11*sw_func_psd_nw_cj} cjswgs = {2.4701E-10*sw_func_psd_nw_cj}
+ mjswgs = 0.70393 pbs = 0.6587 pbsws = 0.7418
+ pbswgs = 1.3925 xrcrg1 = 12 xrcrg2 = 1
+ rbpb = 50 rbpd = 50 rbps = 50
+ rbdb = 50 rbsb = 50 gbmin = 1E-12
+ tnom = 30 ute = 0.949042029246579 wute = -1.061057410227488E-6
+ kt1 = -0.454592552886044 wkt1 = 1.356221220759459E-8 kt1l = 0
+ kt2 = -0.056843931840338 wkt2 = 4.401456148447937E-9 ua1 = 4.482777573077512E-9
+ wua1 = -2.610235795379316E-15 ub1 = -2.617576331055467E-18 wub1 = 1.8660726484721E-24
+ uc1 = -9.810947945401426E-11 wuc1 = 8.767489451919706E-17 at = -7.29161882824356E4
+ wat = 0.071550613908282 prt = 0 njs = 1.2556
+ xtis = 2 tpb = 1.9551E-3 tpbsw = 1.4242E-4
+ tpbswg = 0 tcj = 1.2407E-3 tcjsw = 0
+ tcjswg = 2E-12 tvoff = 0 tvfbsdoff = 0
+ saref = 3E-6 sbref = 3E-6 wlod = 0
+ ku0 = 4.5E-8 kvsat = 0.4 kvth0 = 2.65E-8
+ tku0 = 0 llodku0 = 0 wlodku0 = 1
+ llodvth = 0 wlodvth = 1 lku0 = 0
+ wku0 = 2.5E-7 pku0 = 0 lkvth0 = 0
+ wkvth0 = 2.5E-7 pkvth0 = 0 stk2 = 0
+ lodk2 = 1 steta0 = 0 lodeta0 = 1

.model phighvt_model.34 pmos
+ level = 54 lmin = 4E-6 lmax = 8E-6 wmin = 5.5E-7
+ wmax = 1E-6 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 4.23E-9
+ toxm = 4.23E-9 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 9.999999999999999E22 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {9.364E-9+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {-1.176E-8-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = -5.722E-9 dwb = -1.7864E-8 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = -1.137558506207206 lvth0 = 2.941374104385365E-7
+ wvth0 = 4.618768076374078E-8 pvth0 = -2.704682467283993E-13 k1 = 0.450079833528231
+ lk1 = -7.733553137169382E-8 wk1 = 5.488302073514868E-9 pk1 = 1.167927941716152E-14
+ k2 = 4.380031133136881E-3 lk2 = 9.437184472037713E-8 wk2 = 1.420288687946837E-8
+ pk2 = -7.582556694154958E-14 k3 = -13.778 k3b = 2
+ w0 = 0 lpe0 = 0 lpeb = 0
+ vbm = -3 dvtp0 = 0 dvtp1 = 0
+ dvt0 = 4.05 dvt1 = 0.3 dvt2 = 0.03
+ dvt0w = -4.254 dvt1w = 1.1472E6 dvt2w = -8.96E-3
+ vfbsdoff = 0 u0 = 0.012003564385571 lu0 = -1.54990548390363E-8
+ wu0 = -3.402349130699288E-9 pu0 = 1.900700484465051E-14 ua = -1.178778800465879E-9
+ lua = 1.500460281059728E-15 wua = 3.483430732739124E-16 pua = -7.080837798680863E-22
+ ub = 2.379563275027761E-18 lub = -5.343854514466495E-24 wub = -1.306116799997424E-24
+ pub = 4.745810593006714E-30 uc = -2.813664322697316E-11 luc = -1.485711933843798E-17
+ wuc = -4.190166598543497E-17 puc = 7.186766994893329E-24 ud = 0
+ up = 0 lp = 1 eu = 1.67
+ vsat = 5.090898213320448E5 lvsat = -1.858323915678167 wvsat = -0.236760733107176
+ pvsat = 9.771430500111787E-7 a0 = 1.54887071243518 la0 = -2.028794234372283E-6
+ wa0 = -2.017068903416974E-7 pa0 = 1.29829766212631E-12 ags = 0.394382401244489
+ lags = 7.469506246552395E-9 wags = -1.857404117323052E-7 pags = 2.916017267759595E-13
+ b0 = -1.362408365037191E-7 lb0 = 8.802722061301114E-13 wb0 = 1.336893181176775E-13
+ pb0 = -8.637864682537065E-19 b1 = 1.725418412829142E-10 lb1 = -1.661030823248772E-15
+ wb1 = -1.693104776793678E-16 pb1 = 1.629923037990969E-21 keta = -0.010726212444769
+ lketa = -1.420211753513694E-8 wketa = 9.704539983121466E-9 pketa = 5.797218475857594E-15
+ a1 = 0 a2 = 0.8 rdsw = 531.92
+ rdswmin = 0 rdw = 0 rdwmin = 0
+ rsw = 0 rswmin = 0 prwb = -0.32348
+ prwg = 0.02 wr = 1 voff = -0.223917790287098
+ lvoff = 1.38376588773099E-8 wvoff = 1.785016698387538E-8 pvoff = -6.320343867181331E-14
+ voffl = 0 minv = 0 nfactor = 3.770057354885549
+ lnfactor = -1.259107113961437E-5 wnfactor = -1.589488201406593E-6 pnfactor = 9.71355068258296E-12
+ eta0 = 0.08 etab = -0.07 dsub = 0.56
+ cit = 1E-5 cdsc = 0 cdscb = 0
+ cdscd = 0 pclm = 1.010050518655837 lpclm = -6.97317334223588E-6
+ wpclm = -7.549290952918022E-7 ppclm = 6.05718869465568E-12 pdiblc1 = 0.39
+ pdiblc2 = -3.32150710466008E-3 lpdiblc2 = 2.909911155969636E-8 wpdiblc2 = 1.887807270327501E-9
+ ppdiblc2 = -1.503601375237066E-14 pdiblcb = -0.278209778724115 lpdiblcb = 1.649567048208066E-6
+ wpdiblcb = 2.826886556231788E-8 ppdiblcb = -8.763687848355955E-13 drout = 0.56
+ pscbe1 = 1.731581608270905E9 lpscbe1 = -7.475416601608163E3 wpscbe1 = -494.9232241893004
+ ppscbe1 = 3.971479528769572E-3 pscbe2 = -5.460125114421012E-8 lpscbe2 = 4.207198431929159E-13
+ wpscbe2 = 3.678322795345393E-14 ppscbe2 = -2.353659103636508E-19 pvag = 0
+ delta = 0.01 fprout = 0 pdits = 0
+ pditsl = 0 pditsd = 0 lambda = 0
+ vtl = 0 lc = 5E-9 xn = 3
+ alpha0 = -1.875463985777775E-11 lalpha0 = 9.528302279916774E-16 walpha0 = 1.165306029625213E-16
+ palpha0 = -9.349856234818493E-22 alpha1 = -1.875463985777775E-11 lalpha1 = 9.528302279916774E-16
+ walpha1 = 1.165306029625213E-16 palpha1 = -9.349856234818493E-22 beta0 = 36.00048881786656
+ lbeta0 = -2.074174791607182E-4 wbeta0 = -3.196092443796561E-5 pbeta0 = 2.259639716896619E-10
+ aigbacc = 0.43 bigbacc = 0.054 cigbacc = 0.075
+ nigbacc = 1 aigbinv = 0.35 bigbinv = 0.03
+ cigbinv = 6E-3 eigbinv = 1.1 nigbinv = 3
+ aigc = 0.43 bigc = 0.054 cigc = 0.075
+ aigsd = 0.43 bigsd = 0.054 cigsd = 0.075
+ dlcig = 0 nigc = 1 poxedge = 1
+ pigcd = 1 ntox = 1 toxref = 4.23E-9
+ agidl = 6.887631819229924E-10 lagidl = -2.823026337290628E-15 wagidl = 3.119334232521239E-18
+ pagidl = 8.266882956823185E-22 bgidl = 1E9 cgidl = 300
+ egidl = 3.535580994741011 legidl = -1.382312884396035E-5 wegidl = -1.825227986238046E-6
+ pegidl = 7.343841307188503E-12 noia = 1.2E41 noib = 2E25
+ noic = 0 em = 4.1E7 af = 1
+ ef = 0.88 kf = 0 lintnoi = -6E-8
+ tnoia = 1.5 tnoib = 3.5 ntnoi = 1
+ rnoia = 0.577 rnoib = 0.37 xpart = 0
+ cgso = {5.932020000000001E-11/sw_func_tox_lv_ratio} cgdo = {5.932020000000001E-11/sw_func_tox_lv_ratio} cgbo = {0/sw_func_tox_lv_ratio}
+ ckappas = 0.6 cf = 1.2E-11 clc = 1E-7
+ cle = 0.6 dlc = -2.56E-9 dwc = 0
+ vfbcv = -0.1446893 noff = 4 voffcv = -0.1375
+ acde = 0.552 moin = 14.504 cgsl = {7.513892E-12/sw_func_tox_lv_ratio}
+ cgdl = {7.513892E-12/sw_func_tox_lv_ratio} ijthsrev = 0.1 ijthsfwd = 0.1
+ xjbvs = 1 bvs = 12.8 jss = 2.17E-5
+ jsws = 8.200000000000001E-10 cjs = {7.433E-04*sw_func_psd_nw_cj} mjs = 0.34629
+ mjsws = 0.26859 cjsws = {9.2435E-11*sw_func_psd_nw_cj} cjswgs = {2.4701E-10*sw_func_psd_nw_cj}
+ mjswgs = 0.70393 pbs = 0.6587 pbsws = 0.7418
+ pbswgs = 1.3925 xrcrg1 = 12 xrcrg2 = 1
+ rbpb = 50 rbpd = 50 rbps = 50
+ rbdb = 50 rbsb = 50 gbmin = 1E-12
+ tnom = 30 ute = 1.905709825471143 lute = -7.675843196363717E-6
+ wute = -2.031656743688814E-6 pute = 7.787623164013617E-12 kt1 = -0.397043570155119
+ lkt1 = -4.617454139212331E-7 wkt1 = -8.89701057481929E-9 pkt1 = 1.802020231791534E-13
+ kt1l = 0 kt2 = -0.060056097784704 lkt2 = 2.577287769794022E-8
+ wkt2 = 1.144490489555736E-8 pkt2 = -5.651325189140737E-14 ua1 = 4.745129855035084E-9
+ lua1 = -2.104988781332219E-15 wua1 = -4.096616602673854E-15 pua1 = 1.192600613494387E-20
+ ub1 = -1.6631940506073E-18 lub1 = -7.65750531482148E-24 wub1 = 2.440538724202153E-24
+ pub1 = -4.60924004794159E-30 uc1 = -6.804352381771486E-10 luc1 = 4.672302371630242E-15
+ wuc1 = 6.562616793557346E-16 puc1 = -4.562067439871656E-21 at = -2.252219450770407E5
+ lat = 1.22202828575665 wat = 0.13150297903679 pat = -4.810290006558895E-7
+ prt = 0 njs = 1.2556 xtis = 2
+ tpb = 1.9551E-3 tpbsw = 1.4242E-4 tpbswg = 0
+ tcj = 1.2407E-3 tcjsw = 0 tcjswg = 2E-12
+ tvoff = 0 tvfbsdoff = 0 saref = 3E-6
+ sbref = 3E-6 wlod = 0 ku0 = 4.5E-8
+ kvsat = 0.4 kvth0 = 2.65E-8 tku0 = 0
+ llodku0 = 0 wlodku0 = 1 llodvth = 0
+ wlodvth = 1 lku0 = 0 wku0 = 2.5E-7
+ pku0 = 0 lkvth0 = 0 wkvth0 = 2.5E-7
+ pkvth0 = 0 stk2 = 0 lodk2 = 1
+ steta0 = 0 lodeta0 = 1

.model phighvt_model.35 pmos
+ level = 54 lmin = 2E-6 lmax = 4E-6 wmin = 5.5E-7
+ wmax = 1E-6 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 4.23E-9
+ toxm = 4.23E-9 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 9.999999999999999E22 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {9.364E-9+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {-1.176E-8-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = -5.722E-9 dwb = -1.7864E-8 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = -1.060793334295703 lvth0 = -1.472879405083193E-8
+ wvth0 = -2.408482336564353E-8 pvth0 = 1.227457908626108E-14 k1 = 0.510651898537388
+ lk1 = -3.210484463773401E-7 wk1 = -6.657404868426187E-8 pk1 = 3.016235889380913E-13
+ k2 = -1.627785500581888E-4 lk2 = 1.126499303369061E-7 wk2 = 2.168241727014513E-8
+ pk2 = -1.059196070590453E-13 k3 = -13.778 k3b = 2
+ w0 = 0 lpe0 = 0 lpeb = 0
+ vbm = -3 dvtp0 = 0 dvtp1 = 0
+ dvt0 = 4.05 dvt1 = 0.3 dvt2 = 0.03
+ dvt0w = -4.254 dvt1w = 1.1472E6 dvt2w = -8.96E-3
+ vfbsdoff = 0 u0 = 4.526010905444411E-3 lu0 = 1.458703113932347E-8
+ wu0 = 4.031108260094129E-9 pu0 = -1.090165963635462E-14 ua = -1.637007725358346E-9
+ lua = 3.344153524943065E-15 wua = 8.001723475352403E-16 pua = -2.526027901444024E-21
+ ub = 1.475193156663076E-18 lub = -1.705103255823819E-24 wub = -4.550050157427398E-25
+ pub = 1.321345306822308E-30 uc = -6.886688893537709E-12 luc = -1.003567355981022E-16
+ wuc = -6.743019784163661E-17 puc = 1.099013254889578E-22 ud = 0
+ up = 0 lp = 1 eu = 1.67
+ vsat = 1.748676041509352E4 lvsat = 0.119650831982404 wvsat = 0.03527794476996
+ pvsat = -1.17410011201038E-7 a0 = 0.909593853597943 la0 = 5.433489926965171E-7
+ wa0 = 2.609455674545471E-7 pa0 = -5.631937548660364E-13 ags = 0.406280687599804
+ lags = -4.040348686978327E-8 wags = -2.39392047601169E-7 pags = 5.074701567270507E-13
+ b0 = 1.185319076844274E-7 lb0 = -1.448110255657803E-13 wb0 = -1.163120421173134E-13
+ pb0 = 1.420990046789843E-19 b1 = -2.350626829963079E-9 lb1 = 8.490988788882907E-15
+ wb1 = 2.306604290691531E-15 pb1 = -8.33196955084471E-21 keta = -0.012585924912002
+ lketa = -6.719527228975984E-9 wketa = 1.880536179479715E-8 pketa = -3.082012009985577E-14
+ a1 = 0 a2 = 0.8 rdsw = 531.92
+ rdswmin = 0 rdw = 0 rdwmin = 0
+ rsw = 0 rswmin = 0 prwb = -0.32348
+ prwg = 0.02 wr = 1 voff = -0.247261008105893
+ lvoff = 1.077595626355856E-7 wvoff = 1.322291175671532E-8 pvoff = -4.458558472023027E-14
+ voffl = 0 minv = 0 nfactor = -0.962427210125789
+ lnfactor = 6.450175157400055E-6 wnfactor = 1.717809507340145E-6 pnfactor = -3.593427794513716E-12
+ eta0 = 0.16043492 leta0 = -3.236315093184E-7 etab = -0.140320075185005
+ letab = 2.829342289083728E-7 wetab = 1.463752648169916E-12 petab = -5.88943805496462E-18
+ dsub = 0.860662117397195 ldsub = -1.209720042589963E-6 wdsub = 1.522557806959732E-9
+ pdsub = -6.126041787458619E-15 cit = 1E-5 cdsc = 0
+ cdscb = 0 cdscd = 0 pclm = -1.927790694004172
+ lpclm = 4.847289533725918E-6 wpclm = 1.34612687090321E-6 ppclm = -2.396452006449276E-12
+ pdiblc1 = 0.39 pdiblc2 = 7.445949838902158E-3 lpdiblc2 = -1.422396680186518E-8
+ wpdiblc2 = -3.733464399179453E-9 ppdiblc2 = 7.581285235323954E-15 pdiblcb = 0.290386219658008
+ lpdiblcb = -6.381903232023717E-7 wpdiblcb = -3.813142194341491E-7 ppdiblcb = 7.715969493093893E-13
+ drout = 0.56 pscbe1 = -1.046470234268693E9 lpscbe1 = 3.70213054788676E3
+ wpscbe1 = 980.9779343003969 ppscbe1 = -1.966838300436895E-3 pscbe2 = 9.11908289469206E-8
+ lpscbe2 = -1.658775068953502E-13 wpscbe2 = -4.381843819431823E-14 ppscbe2 = 8.893650541523334E-20
+ pvag = 0 delta = 0.01 fprout = 0
+ pdits = 0 pditsl = 0 pditsd = 0
+ lambda = 0 vtl = 0 lc = 5E-9
+ xn = 3 alpha0 = 3.375092797155556E-10 lalpha0 = -4.806047776900211E-16
+ walpha0 = -2.330612059250427E-16 palpha0 = 4.716040114134424E-22 alpha1 = 3.375092797155556E-10
+ lalpha1 = -4.806047776900211E-16 walpha1 = -2.330612059250427E-16 palpha1 = 4.716040114134424E-22
+ beta0 = -39.58263445201758 lbeta0 = 9.669272897812598E-5 wbeta0 = 5.010004439395806E-5
+ pbeta0 = -1.042099776249596E-10 aigbacc = 0.43 bigbacc = 0.054
+ cigbacc = 0.075 nigbacc = 1 aigbinv = 0.35
+ bigbinv = 0.03 cigbinv = 6E-3 eigbinv = 1.1
+ nigbinv = 3 aigc = 0.43 bigc = 0.054
+ cigc = 0.075 aigsd = 0.43 bigsd = 0.054
+ cigsd = 0.075 dlcig = 0 nigc = 1
+ poxedge = 1 pigcd = 1 ntox = 1
+ toxref = 4.23E-9 agidl = 6.753314031271871E-10 lagidl = -2.768983306670129E-15
+ wagidl = -3.97829043613243E-16 pagidl = 2.439912112912308E-21 bgidl = 1E9
+ cgidl = 300 egidl = 0.1 noia = 1.2E41
+ noib = 2E25 noic = 0 em = 4.1E7
+ af = 1 ef = 0.88 kf = 0
+ lintnoi = -6E-8 tnoia = 1.5 tnoib = 3.5
+ ntnoi = 1 rnoia = 0.577 rnoib = 0.37
+ xpart = 0 cgso = {5.932020000000001E-11/sw_func_tox_lv_ratio} cgdo = {5.932020000000001E-11/sw_func_tox_lv_ratio}
+ cgbo = {0/sw_func_tox_lv_ratio} ckappas = 0.6 cf = 1.2E-11
+ clc = 1E-7 cle = 0.6 dlc = -2.56E-9
+ dwc = 0 vfbcv = -0.1446893 noff = 4
+ voffcv = -0.1375 acde = 0.552 moin = 14.504
+ cgsl = {7.513892E-12/sw_func_tox_lv_ratio} cgdl = {7.513892E-12/sw_func_tox_lv_ratio} ijthsrev = 0.1
+ ijthsfwd = 0.1 xjbvs = 1 bvs = 12.8
+ jss = 2.17E-5 jsws = 8.200000000000001E-10 cjs = {7.433E-04*sw_func_psd_nw_cj}
+ mjs = 0.34629 mjsws = 0.26859 cjsws = {9.2435E-11*sw_func_psd_nw_cj}
+ cjswgs = {2.4701E-10*sw_func_psd_nw_cj} mjswgs = 0.70393 pbs = 0.6587
+ pbsws = 0.7418 pbswgs = 1.3925 xrcrg1 = 12
+ xrcrg2 = 1 rbpb = 50 rbpd = 50
+ rbps = 50 rbdb = 50 rbsb = 50
+ gbmin = 1E-12 tnom = 30 ute = -0.181366933583177
+ lute = 7.215518852265183E-7 wute = 4.77186835741277E-8 pute = -5.787854550873751E-13
+ kt1 = -0.536023042394866 lkt1 = 9.744127222483207E-8 wkt1 = 5.338986809937156E-8
+ pkt1 = -7.041047890402694E-14 kt1l = 0 kt2 = -0.0568331694892
+ lkt2 = 1.280536124241582E-8 wkt2 = -3.388482498591481E-9 pkt2 = 3.16917895669836E-15
+ ua1 = 3.83925953552953E-9 lua1 = 1.539798566604771E-15 wua1 = -5.059295475678443E-16
+ pua1 = -2.521195045016262E-21 ub1 = -3.94914493554688E-18 lub1 = 1.540063789750625E-24
+ wub1 = 1.086093264435495E-24 pub1 = 8.403983483387532E-31 uc1 = 1.07521107912521E-9
+ luc1 = -2.391575698962144E-15 wuc1 = -1.037230053368476E-15 puc1 = 2.251730416578861E-21
+ at = 3.103412572149756E4 lat = 0.190976859777315 wat = 0.069926351494155
+ pat = -2.332742082055451E-7 prt = 0 njs = 1.2556
+ xtis = 2 tpb = 1.9551E-3 tpbsw = 1.4242E-4
+ tpbswg = 0 tcj = 1.2407E-3 tcjsw = 0
+ tcjswg = 2E-12 tvoff = 0 tvfbsdoff = 0
+ saref = 3E-6 sbref = 3E-6 wlod = 0
+ ku0 = 4.5E-8 kvsat = 0.4 kvth0 = 2.65E-8
+ tku0 = 0 llodku0 = 0 wlodku0 = 1
+ llodvth = 0 wlodvth = 1 lku0 = 0
+ wku0 = 2.5E-7 pku0 = 0 lkvth0 = 0
+ wkvth0 = 2.5E-7 pkvth0 = 0 stk2 = 0
+ lodk2 = 1 steta0 = 0 lodeta0 = 1

.model phighvt_model.36 pmos
+ level = 54 lmin = 1E-6 lmax = 2E-6 wmin = 5.5E-7
+ wmax = 1E-6 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 4.23E-9
+ toxm = 4.23E-9 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 9.999999999999999E22 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {9.364E-9+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {-1.176E-8-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = -5.722E-9 dwb = -1.7864E-8 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = -1.082101734615847 lvth0 = 2.838918016498516E-8
+ wvth0 = -1.912836810400784E-8 pvth0 = 2.245092735236027E-15 k1 = 0.174070096422376
+ lk1 = 3.600315618384294E-7 wk1 = 1.765922364402255E-7 pk1 = -1.904282523370114E-13
+ k2 = 0.124886767335908 lk2 = -1.40390326754265E-7 wk2 = -6.7814989371245E-8
+ pk2 = 7.51801852279404E-14 k3 = -13.778 k3b = 2
+ w0 = 0 lpe0 = 0 lpeb = 0
+ vbm = -3 dvtp0 = 0 dvtp1 = 0
+ dvt0 = 4.05 dvt1 = 0.3 dvt2 = 0.03
+ dvt0w = -4.254 dvt1w = 1.1472E6 dvt2w = -8.96E-3
+ vfbsdoff = 0 u0 = 0.01373635979908 lu0 = -4.050294053926842E-9
+ wu0 = -1.209842158863068E-9 pu0 = -2.964916445863532E-16 ua = 4.49186547430914E-10
+ lua = -8.773023099314574E-16 wua = -4.149370574601541E-16 pua = -6.722971824774386E-23
+ ub = 4.615059858763586E-19 lub = 3.461130080065193E-25 wub = 1.336366821984552E-25
+ pub = 1.302170582043417E-31 uc = -2.24896572351309E-11 luc = -6.878381709952153E-17
+ wuc = -5.161695680377568E-17 puc = 7.790291598402543E-23 ud = 0
+ up = 0 lp = 1 eu = 1.67
+ vsat = 1.118973919899224E5 lvsat = -0.071390969221893 wvsat = -0.051280203004084
+ pvsat = 5.774213198269547E-8 a0 = 1.764126054292167 la0 = -1.185814006052258E-6
+ wa0 = -3.895220023122443E-7 pa0 = 7.530403819084614E-13 ags = 0.090452822727839
+ lags = 5.986805142559346E-7 wags = 8.347126665104783E-8 pags = -1.458502169285952E-13
+ b0 = -1.83372838589497E-8 lb0 = 1.321465209060742E-13 wb0 = 1.799386320683928E-14
+ pb0 = -1.296716808625452E-19 b1 = 3.58374019752687E-9 lb1 = -3.517321578583553E-15
+ wb1 = -3.516623911107587E-15 pb1 = 3.45144918005984E-21 keta = -2.874558076547403E-3
+ lketa = -2.637067224785452E-8 wketa = -7.776369433653534E-9 pketa = 2.296854467553876E-14
+ a1 = 0 a2 = 0.353621547804445 la2 = 9.032557255867503E-7
+ wa2 = 2.371483730548372E-7 pa2 = -4.798744758439241E-13 rdsw = 531.92
+ rdswmin = 0 rdw = 0 rdwmin = 0
+ rsw = 0 rswmin = 0 prwb = -0.32348
+ prwg = 0.02 wr = 1 voff = -0.198557651033484
+ lvoff = 9.207345532426235E-9 wvoff = -3.550872942536977E-9 pvoff = -1.064349590559926E-14
+ voffl = 0 minv = 0 nfactor = 2.338790690392377
+ lnfactor = -2.299052886564636E-7 wnfactor = 8.996458164885985E-8 pnfactor = -2.994510304788878E-13
+ eta0 = 0.102097870464 leta0 = -2.055853228413134E-7 weta0 = -3.201503036240302E-7
+ peta0 = 6.478305423892977E-13 etab = 1.840771095127327 letab = -3.725843376042038E-6
+ wetab = -9.778095974335504E-7 petab = 1.978614349093441E-12 dsub = -0.887662102627327
+ ldsub = 2.328048983114059E-6 wdsub = 6.097207513374206E-7 pdsub = -1.236827250360217E-12
+ cit = 1E-5 cdsc = 0 cdscb = 0
+ cdscd = 0 pclm = -0.09383543134625 lpclm = 1.136244380632362E-6
+ wpclm = 5.38578500345439E-7 ppclm = -7.62361727658215E-13 pdiblc1 = 1.166553757405921
+ lpdiblc1 = -1.57137205918603E-6 wpdiblc1 = -4.094830760157832E-7 ppdiblc1 = 8.285971939794577E-13
+ pdiblc2 = 4.029480161501114E-4 lpdiblc2 = 2.768824651003788E-11 wpdiblc2 = 2.65453542963478E-11
+ ppdiblc2 = -2.716970102939789E-17 pdiblcb = -0.266674452195555 lpdiblcb = 4.890330875067505E-7
+ wpdiblcb = 2.371483730548372E-7 ppdiblcb = -4.798744758439242E-13 drout = -0.208917453087914
+ ldrout = 1.555919844672455E-6 wdrout = 3.126024993528834E-7 pdrout = -6.325574094905466E-13
+ pscbe1 = 7.963329793382609E8 lpscbe1 = -26.818610911182493 wpscbe1 = 1.948185401003484
+ ppscbe1 = 1.424797705600575E-5 pscbe2 = 9.248348370310011E-9 lpscbe2 = -6.525859896721196E-17
+ wpscbe2 = 2.768872318393766E-16 ppscbe2 = -2.912674911050781E-22 pvag = 0
+ delta = 0.01 fprout = 0 pdits = 0
+ pditsl = 0 pditsd = 0 lambda = 0
+ vtl = 0 lc = 5E-9 xn = 3
+ alpha0 = 1E-10 alpha1 = 1E-10 beta0 = 7.301555985893016
+ lbeta0 = 1.821631943205164E-6 wbeta0 = -1.412288272152907E-6 pbeta0 = 2.625777156922797E-14
+ aigbacc = 0.43 bigbacc = 0.054 cigbacc = 0.075
+ nigbacc = 1 aigbinv = 0.35 bigbinv = 0.03
+ cigbinv = 6E-3 eigbinv = 1.1 nigbinv = 3
+ aigc = 0.43 bigc = 0.054 cigc = 0.075
+ aigsd = 0.43 bigsd = 0.054 cigsd = 0.075
+ dlcig = 0 nigc = 1 poxedge = 1
+ pigcd = 1 ntox = 1 toxref = 4.23E-9
+ agidl = -1.045105721667239E-9 lagidl = 7.123556240938883E-16 wagidl = 7.739904384692557E-16
+ pagidl = 6.871195452873031E-23 bgidl = 1E9 cgidl = 300
+ egidl = 0.1 noia = 1.2E41 noib = 2E25
+ noic = 0 em = 4.1E7 af = 1
+ ef = 0.88 kf = 0 lintnoi = -6E-8
+ tnoia = 1.5 tnoib = 3.5 ntnoi = 1
+ rnoia = 0.577 rnoib = 0.37 xpart = 0
+ cgso = {5.932020000000001E-11/sw_func_tox_lv_ratio} cgdo = {5.932020000000001E-11/sw_func_tox_lv_ratio} cgbo = {0/sw_func_tox_lv_ratio}
+ ckappas = 0.6 cf = 1.2E-11 clc = 1E-7
+ cle = 0.6 dlc = -2.56E-9 dwc = 0
+ vfbcv = -0.1446893 noff = 4 voffcv = -0.1375
+ acde = 0.552 moin = 14.504 cgsl = {7.513892E-12/sw_func_tox_lv_ratio}
+ cgdl = {7.513892E-12/sw_func_tox_lv_ratio} ijthsrev = 0.1 ijthsfwd = 0.1
+ xjbvs = 1 bvs = 12.8 jss = 2.17E-5
+ jsws = 8.200000000000001E-10 cjs = {7.433E-04*sw_func_psd_nw_cj} mjs = 0.34629
+ mjsws = 0.26859 cjsws = {9.2435E-11*sw_func_psd_nw_cj} cjswgs = {2.4701E-10*sw_func_psd_nw_cj}
+ mjswgs = 0.70393 pbs = 0.6587 pbsws = 0.7418
+ pbswgs = 1.3925 xrcrg1 = 12 xrcrg2 = 1
+ rbpb = 50 rbpd = 50 rbps = 50
+ rbdb = 50 rbsb = 50 gbmin = 1E-12
+ tnom = 30 ute = 1.427364786278289 lute = -2.533748924547554E-6
+ wute = -4.822257445014563E-7 pute = 4.935676940121305E-13 kt1 = -0.496879731837227
+ lkt1 = 1.823400044523829E-8 wkt1 = 3.762498699241338E-8 pkt1 = -3.850992668647494E-14
+ kt1l = 0 kt2 = -0.052496400945251 lkt2 = 4.029823358363146E-9
+ wkt2 = -3.687483148851473E-9 pkt2 = 3.774212752512459E-15 ua1 = 9.749144113784283E-9
+ lua1 = -1.041897107518529E-14 wua1 = -3.544953603110746E-15 pua1 = 3.62833091185591E-21
+ ub1 = -7.415378118802309E-18 lub1 = 8.55405596073165E-24 wub1 = 3.085559465400232E-24
+ pub1 = -3.205561498637412E-30 uc1 = -2.843572878833394E-10 luc1 = 3.595380830469955E-16
+ wuc1 = 1.528746589866824E-16 puc1 = -1.564702709660492E-22 at = 1.784769320521422E5
+ lat = -0.107376607688871 wat = -0.079919418777351 pat = 6.994170485425195E-8
+ prt = 0 njs = 1.2556 xtis = 2
+ tpb = 1.9551E-3 tpbsw = 1.4242E-4 tpbswg = 0
+ tcj = 1.2407E-3 tcjsw = 0 tcjswg = 2E-12
+ tvoff = 0 tvfbsdoff = 0 saref = 3E-6
+ sbref = 3E-6 wlod = 0 ku0 = 4.5E-8
+ kvsat = 0.4 kvth0 = 2.65E-8 tku0 = 0
+ llodku0 = 0 wlodku0 = 1 llodvth = 0
+ wlodvth = 1 lku0 = 0 wku0 = 2.5E-7
+ pku0 = 0 lkvth0 = 0 wkvth0 = 2.5E-7
+ pkvth0 = 0 stk2 = 0 lodk2 = 1
+ steta0 = 0 lodeta0 = 1

.model phighvt_model.37 pmos
+ level = 54 lmin = 5E-7 lmax = 1E-6 wmin = 5.5E-7
+ wmax = 1E-6 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 4.23E-9
+ toxm = 4.23E-9 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 9.999999999999999E22 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {9.364E-9+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {-1.176E-8-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = -5.722E-9 dwb = -1.7864E-8 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = -1.079905341678665 lvth0 = 2.614112806592022E-8
+ wvth0 = -1.287304939682645E-8 pvth0 = -4.157351067938271E-15 k1 = 0.435848320418169
+ lk1 = 9.209631401425581E-8 wk1 = 7.899267974405321E-8 pk1 = -9.053315406734516E-14
+ k2 = 0.015634502598809 lk2 = -2.856844875054853E-8 wk2 = -2.701640883669354E-8
+ pk2 = 3.34220220792163E-14 k3 = -13.778 k3b = 2
+ w0 = 0 lpe0 = 0 lpeb = 0
+ vbm = -3 dvtp0 = 0 dvtp1 = 0
+ dvt0 = 4.05 dvt1 = 0.3 dvt2 = 0.03
+ dvt0w = -4.254 dvt1w = 1.1472E6 dvt2w = -8.96E-3
+ vfbsdoff = 0 u0 = 0.015379746399101 lu0 = -5.732333106780293E-9
+ wu0 = -5.380117649707635E-9 pu0 = 3.971868725802877E-15 ua = 1.002116194442195E-9
+ lua = -1.443236862240443E-15 wua = -1.518037765427145E-15 pua = 1.061815918370631E-21
+ ub = -6.542702204415059E-20 lub = 8.854394802733187E-25 wub = 9.097308059325721E-25
+ pub = -6.641307993200016E-31 uc = -1.754737760018781E-10 luc = 8.779848814061951E-17
+ wuc = 7.270962589812021E-17 puc = -4.934782794301904E-23 ud = 0
+ up = 0 lp = 1 eu = 1.67
+ vsat = -1.941565325115219E4 lvsat = 0.063010558843251 wvsat = 0.013115925978173
+ pvsat = -8.16859395322391E-9 a0 = 0.981163780708417 la0 = -3.844364597938182E-7
+ wa0 = 2.261742330729183E-7 pa0 = 1.228629710670399E-13 ags = 0.073721574748666
+ lags = 6.158052811875785E-7 wags = -1.208314121718294E-7 pags = 6.325766090019612E-14
+ b0 = 2.26755888261524E-7 lb0 = -1.18711242622673E-13 wb0 = -2.225092039861621E-13
+ pb0 = 1.164880184708356E-19 b1 = 3.014163767782971E-10 lb1 = -1.57797501570974E-16
+ wb1 = -2.957714508739931E-16 pb1 = 1.548422699615528E-22 keta = -0.026319107411297
+ lketa = -2.374707112751891E-9 wketa = 3.706965887862021E-8 pketa = -2.293226222263966E-14
+ a1 = 0 a2 = 0.878209436819513 la2 = 3.66329529422048E-7
+ wa2 = 1.296917371037316E-7 pa2 = -3.698904598152486E-13 rdsw = 531.92
+ rdswmin = 0 rdw = 0 rdwmin = 0
+ rsw = 0 rswmin = 0 prwb = -0.32348
+ prwg = 0.02 wr = 1 voff = -0.164296594809518
+ lvoff = -2.585953073392799E-8 wvoff = -3.418657786593704E-8 pvoff = 2.071276079759917E-14
+ voffl = 0 minv = 0 nfactor = 3.289986643847975
+ lnfactor = -1.203473370937337E-6 wnfactor = -1.463741930256526E-6 pnfactor = 1.290798658586512E-12
+ eta0 = -1.310830534005536 leta0 = 1.240575157701346E-6 weta0 = 1.22475476034708E-6
+ peta0 = -9.334106886864128E-13 etab = -3.68336384072103 letab = 1.928219213497472E-6
+ wetab = 1.956068209675912E-6 petab = -1.024268264039235E-12 dsub = 3.475712617269356
+ ldsub = -2.137952310194594E-6 wdsub = -2.120052719413125E-6 pdsub = 1.557150492422382E-12
+ cit = 1E-5 cdsc = 0 cdscb = 0
+ cdscd = 0 pclm = 2.5514651226346 lpclm = -1.571273642378117E-6
+ wpclm = -9.130806931981467E-7 ppclm = 7.234404901175156E-13 pdiblc1 = -0.693505593182428
+ lpdiblc1 = 3.324358873281566E-7 wpdiblc1 = 7.475550025372399E-7 ppdiblc1 = -3.556544201811323E-13
+ pdiblc2 = 1.781990405424078E-3 lpdiblc2 = -1.383789219759651E-9 wpdiblc2 = -9.261113879594762E-10
+ ppdiblc2 = 9.47893527804283E-16 pdiblcb = 0.198629948595477 lpdiblcb = 1.278472720911286E-8
+ wpdiblcb = -2.250627300502164E-7 ppdiblcb = -6.792167593839809E-15 drout = 1.033870106655471
+ ldrout = 2.839019215239057E-7 wdrout = -3.323578729802784E-8 pdrout = -2.78585006337606E-13
+ pscbe1 = -7.911652494585776E7 lpscbe1 = 869.2214657136982 wpscbe1 = 835.1377387576744
+ ppscbe1 = -8.385381945956139E-4 pscbe2 = 9.413844816524973E-8 lpscbe2 = -8.695197354108386E-14
+ wpscbe2 = -8.352607729195474E-14 ppscbe2 = 8.548274275828866E-20 pvag = 0
+ delta = 0.01 fprout = 0 pdits = 0
+ pditsl = 0 pditsd = 0 lambda = 0
+ vtl = 0 lc = 5E-9 xn = 3
+ alpha0 = 1E-10 alpha1 = 1E-10 beta0 = 9.04406571758671
+ lbeta0 = 3.81383826220345E-8 wbeta0 = -2.463131513924702E-6 pbeta0 = 1.101816846387495E-12
+ aigbacc = 0.43 bigbacc = 0.054 cigbacc = 0.075
+ nigbacc = 1 aigbinv = 0.35 bigbinv = 0.03
+ cigbinv = 6E-3 eigbinv = 1.1 nigbinv = 3
+ aigc = 0.43 bigc = 0.054 cigc = 0.075
+ aigsd = 0.43 bigsd = 0.054 cigsd = 0.075
+ dlcig = 0 nigc = 1 poxedge = 1
+ pigcd = 1 ntox = 1 toxref = 4.23E-9
+ agidl = -2.524716707422489E-11 lagidl = -3.314900037031535E-16 wagidl = 8.474575843039875E-16
+ pagidl = -6.483138576034395E-24 bgidl = 1E9 cgidl = 300
+ egidl = 0.1 noia = 1.2E41 noib = 2E25
+ noic = 0 em = 4.1E7 af = 1
+ ef = 0.88 kf = 0 lintnoi = -6E-8
+ tnoia = 1.5 tnoib = 3.5 ntnoi = 1
+ rnoia = 0.577 rnoib = 0.37 xpart = 0
+ cgso = {5.932020000000001E-11/sw_func_tox_lv_ratio} cgdo = {5.932020000000001E-11/sw_func_tox_lv_ratio} cgbo = {0/sw_func_tox_lv_ratio}
+ ckappas = 0.6 cf = 1.2E-11 clc = 1E-7
+ cle = 0.6 dlc = -2.56E-9 dwc = 0
+ vfbcv = -0.1446893 noff = 4 voffcv = -0.1375
+ acde = 0.552 moin = 14.504 cgsl = {7.513892E-12/sw_func_tox_lv_ratio}
+ cgdl = {7.513892E-12/sw_func_tox_lv_ratio} ijthsrev = 0.1 ijthsfwd = 0.1
+ xjbvs = 1 bvs = 12.8 jss = 2.17E-5
+ jsws = 8.200000000000001E-10 cjs = {7.433E-04*sw_func_psd_nw_cj} mjs = 0.34629
+ mjsws = 0.26859 cjsws = {9.2435E-11*sw_func_psd_nw_cj} cjswgs = {2.4701E-10*sw_func_psd_nw_cj}
+ mjswgs = 0.70393 pbs = 0.6587 pbsws = 0.7418
+ pbswgs = 1.3925 xrcrg1 = 12 xrcrg2 = 1
+ rbpb = 50 rbpd = 50 rbps = 50
+ rbdb = 50 rbsb = 50 gbmin = 1E-12
+ tnom = 30 ute = -1.98724265509632 lute = 9.611700838481853E-7
+ wute = 4.858023532788621E-8 pute = -4.972284246279809E-14 kt1 = -0.350297441769273
+ lkt1 = -1.31795905085114E-7 wkt1 = -6.573190892429869E-8 pkt1 = 6.727792342219819E-14
+ kt1l = 0 kt2 = -0.098427233417661 lkt2 = 5.104094901052454E-8
+ wkt2 = 3.260394869858317E-8 pkt2 = -3.337079357197384E-14 ua1 = -4.681920939519361E-9
+ lua1 = 4.351512628172055E-15 wua1 = 1.092782372207061E-15 pua1 = -1.118484613601371E-21
+ ub1 = 6.425258025410091E-18 lub1 = -5.612111945592624E-24 wub1 = -2.001873151296585E-24
+ pub1 = 2.001527533204113E-30 uc1 = 4.997061899652296E-10 luc1 = -4.429665678005717E-16
+ wuc1 = -1.552396279025772E-16 puc1 = 1.588908639508458E-22 at = 1.693683377112221E5
+ lat = -0.098053779209052 wat = -0.078188989323962 pat = 6.817057570011949E-8
+ prt = 0 njs = 1.2556 xtis = 2
+ tpb = 1.9551E-3 tpbsw = 1.4242E-4 tpbswg = 0
+ tcj = 1.2407E-3 tcjsw = 0 tcjswg = 2E-12
+ tvoff = 0 tvfbsdoff = 0 saref = 2.75E-6
+ sbref = 2.74E-6 wlod = 0 ku0 = 4.5E-8
+ kvsat = 0.4 kvth0 = 2.65E-8 tku0 = 0
+ llodku0 = 0 wlodku0 = 1 llodvth = 0
+ wlodvth = 1 lku0 = 0 wku0 = 2.5E-7
+ pku0 = 0 lkvth0 = 0 wkvth0 = 2.5E-7
+ pkvth0 = 0 stk2 = 0 lodk2 = 1
+ steta0 = 0 lodeta0 = 1

.model phighvt_model.38 pmos
+ level = 54 lmin = 2.5E-7 lmax = 5E-7 wmin = 5.5E-7
+ wmax = 1E-6 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 4.23E-9
+ toxm = 4.23E-9 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 9.999999999999999E22 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {9.364E-9+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {-1.176E-8-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = -5.722E-9 dwb = -1.7864E-8 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = -1.03524712017109 lvth0 = 2.761655942274289E-9
+ wvth0 = -1.795817539804715E-8 pvth0 = -1.49518590377921E-15 k1 = 1.101520473011948
+ lk1 = -2.563963713116396E-7 wk1 = -5.963386791378238E-7 pk1 = 2.630163189344951E-13
+ k2 = -0.231660948433154 lk2 = 1.008956657737044E-7 wk2 = 2.262643022708277E-7
+ pk2 = -9.917549579979319E-14 k3 = -13.778 k3b = 2
+ w0 = 0 lpe0 = 0 lpeb = 0
+ vbm = -3 dvtp0 = 0 dvtp1 = 0
+ dvt0 = 4.05 dvt1 = 0.3 dvt2 = 0.03
+ dvt0w = -4.254 dvt1w = 1.1472E6 dvt2w = -8.96E-3
+ vfbsdoff = 0 u0 = -2.059638258217988E-3 lu0 = 3.397533549019534E-9
+ wu0 = 9.304689475433255E-9 pu0 = -3.715921500350881E-15 ua = -4.143556476379676E-9
+ lua = 1.250625694388222E-15 wua = 2.857711704737232E-15 pua = -1.228976444249824E-21
+ ub = 3.449625175676524E-18 lub = -9.547606462774086E-25 wub = -2.142907204534501E-24
+ pub = 9.339862519197207E-31 uc = -1.604250209312335E-11 luc = 4.333027623908246E-18
+ wuc = -4.539823037628088E-17 puc = 1.248399697375541E-23 ud = 0
+ up = 0 lp = 1 eu = 1.67
+ vsat = 9.076352145066609E4 lvsat = 5.32955730335547E-3 wvsat = 8.16351815102717E-3
+ pvsat = -5.575909407556478E-9 a0 = 0.60839865516945 la0 = -1.892864612716584E-7
+ wa0 = 2.385372888322494E-7 pa0 = 1.163906641159148E-13 ags = 0.587714214743609
+ lags = 3.46719854297426E-7 wags = 3.518538937047336E-7 pags = -1.842025504323021E-13
+ b0 = 0 b1 = 0 keta = -0.021588310417523
+ lketa = -4.851373954932452E-9 wketa = -2.055785060333919E-8 pketa = 7.236891541355724E-15
+ a1 = 0 a2 = 1.980232394430791 la2 = -2.106015293466085E-7
+ wa2 = -7.675207233768681E-7 pa2 = 9.981820749555496E-14 rdsw = 531.92
+ rdswmin = 0 rdw = 0 rdwmin = 0
+ rsw = 0 rswmin = 0 prwb = -0.32348
+ prwg = 0.02 wr = 1 voff = -0.267598246133347
+ lvoff = 2.822094976712292E-8 wvoff = 6.752505444291059E-8 pvoff = -3.253531294872874E-14
+ voffl = 0 minv = 0 nfactor = -1.246120958667721
+ lnfactor = 1.17126968113168E-6 wnfactor = 2.745244141672964E-6 pnfactor = -9.12689729790014E-13
+ eta0 = 1.681217426155071 leta0 = -3.258217904019349E-7 weta0 = -1.168908306198039E-6
+ peta0 = 3.197197999112875E-13 etab = -3.748595872064326E-4 letab = 1.008220942927034E-10
+ wetab = -9.097396388067696E-10 petab = 2.488319860064276E-16 dsub = -2.360273838100551
+ ldsub = 9.173033189206593E-7 wdsub = 1.98160440772951E-6 pdsub = -5.901490467793306E-13
+ cit = 1E-5 cdsc = 0 cdscb = 0
+ cdscd = 0 pclm = -1.397847660401928 lpclm = 4.962705857971656E-7
+ wpclm = 7.433128735200657E-7 ppclm = -1.437146699308028E-13 pdiblc1 = -0.855262744423176
+ lpdiblc1 = 4.171189911457136E-7 wpdiblc1 = 4.229709675010388E-7 ppdiblc1 = -1.857281861589803E-13
+ pdiblc2 = -6.875092577055518E-3 lpdiblc2 = 3.148366863228067E-9 wpdiblc2 = -3.041142885086556E-9
+ ppdiblc2 = 2.055154817180252E-15 pdiblcb = 0.692944736668947 lpdiblcb = -2.4599895064311E-7
+ wpdiblcb = -4.876783361395849E-7 ppdiblcb = 1.306923545060664E-13 drout = 3.423050622787258
+ ldrout = -9.668818622814067E-7 wdrout = -1.829137546697708E-6 pdrout = 6.616054827433148E-13
+ pscbe1 = 2.435973974722896E9 lpscbe1 = -447.47871267288724 wpscbe1 = -1.605304373691766E3
+ ppscbe1 = 4.390820601139168E-4 pscbe2 = -1.604806105225941E-7 lpscbe2 = 4.634619606317613E-14
+ wpscbe2 = 1.668145957065018E-13 ppscbe2 = -4.557560636986332E-20 pvag = 0
+ delta = 0.01 fprout = 0 pdits = 0
+ pditsl = 0 pditsd = 0 lambda = 0
+ vtl = 0 lc = 5E-9 xn = 3
+ alpha0 = 1E-10 alpha1 = 1E-10 beta0 = 9.458251821320086
+ lbeta0 = -1.786963264044629E-7 wbeta0 = -9.136430128259946E-7 pbeta0 = 2.906286262923004E-13
+ aigbacc = 0.43 bigbacc = 0.054 cigbacc = 0.075
+ nigbacc = 1 aigbinv = 0.35 bigbinv = 0.03
+ cigbinv = 6E-3 eigbinv = 1.1 nigbinv = 3
+ aigc = 0.43 bigc = 0.054 cigc = 0.075
+ aigsd = 0.43 bigsd = 0.054 cigsd = 0.075
+ dlcig = 0 nigc = 1 poxedge = 1
+ pigcd = 1 ntox = 1 toxref = 4.23E-9
+ agidl = 6.504729004788944E-10 lagidl = -6.852429734685625E-16 wagidl = -3.49945308784491E-16
+ pagidl = 6.203812240136458E-22 bgidl = 3.788257957238561E8 lbgidl = 325.1971194226468
+ wbgidl = 330.0124618541956 pbgidl = -1.727681240299084E-4 cgidl = 300
+ egidl = 0.1 noia = 1.2E41 noib = 2E25
+ noic = 0 em = 4.1E7 af = 1
+ ef = 0.88 kf = 0 lintnoi = -6E-8
+ tnoia = 1.5 tnoib = 3.5 ntnoi = 1
+ rnoia = 0.577 rnoib = 0.37 xpart = 0
+ cgso = {5.932020000000001E-11/sw_func_tox_lv_ratio} cgdo = {5.932020000000001E-11/sw_func_tox_lv_ratio} cgbo = {0/sw_func_tox_lv_ratio}
+ ckappas = 0.6 cf = 1.2E-11 clc = 1E-7
+ cle = 0.6 dlc = -2.56E-9 dwc = 0
+ vfbcv = -0.1446893 noff = 4 voffcv = -0.1375
+ acde = 0.552 moin = 14.504 cgsl = {7.513892E-12/sw_func_tox_lv_ratio}
+ cgdl = {7.513892E-12/sw_func_tox_lv_ratio} ijthsrev = 0.1 ijthsfwd = 0.1
+ xjbvs = 1 bvs = 12.8 jss = 2.17E-5
+ jsws = 8.200000000000001E-10 cjs = {7.433E-04*sw_func_psd_nw_cj} mjs = 0.34629
+ mjsws = 0.26859 cjsws = {9.2435E-11*sw_func_psd_nw_cj} cjswgs = {2.4701E-10*sw_func_psd_nw_cj}
+ mjswgs = 0.70393 pbs = 0.6587 pbsws = 0.7418
+ pbswgs = 1.3925 xrcrg1 = 12 xrcrg2 = 1
+ rbpb = 50 rbpd = 50 rbps = 50
+ rbdb = 50 rbsb = 50 gbmin = 1E-12
+ tnom = 30 ute = 1.799713312966828 lute = -1.021377104552234E-6
+ wute = -1.246291053178258E-6 pute = 6.281681744959383E-13 kt1 = -0.80278303459779
+ lkt1 = 1.050893524724714E-7 wkt1 = 2.375704801354996E-7 pkt1 = -9.150694329838738E-14
+ kt1l = 0 kt2 = 0.069774651468274 lkt2 = -3.701610176495997E-8
+ wkt2 = -7.870734239749198E-8 pkt2 = 2.490289354264341E-14 ua1 = 7.287754322031166E-9
+ lua1 = -1.914851764754876E-15 wua1 = -2.189255648664587E-15 pua1 = 5.997279310853542E-22
+ ub1 = -8.507872304383767E-18 lub1 = 2.205680444661055E-24 wub1 = 3.524335887408637E-24
+ pub1 = -8.915534227388443E-31 uc1 = -5.81762208671821E-10 luc1 = 1.232037682538969E-16
+ wuc1 = 2.807692060724726E-16 puc1 = -6.936848081177224E-23 at = -1.125268940850962E5
+ lat = 0.049524012540956 wat = 0.105166587006317 pat = -2.781973562030807E-8
+ prt = 0 njs = 1.2556 xtis = 2
+ tpb = 1.9551E-3 tpbsw = 1.4242E-4 tpbswg = 0
+ tcj = 1.2407E-3 tcjsw = 0 tcjswg = 2E-12
+ tvoff = 0 tvfbsdoff = 0 saref = 1.75E-6
+ sbref = 1.74E-6 wlod = 0 ku0 = 4.5E-8
+ kvsat = 0.4 kvth0 = 2.65E-8 tku0 = 0
+ llodku0 = 0 wlodku0 = 1 llodvth = 0
+ wlodvth = 1 lku0 = 0 wku0 = 2.5E-7
+ pku0 = 0 lkvth0 = 0 wkvth0 = 2.5E-7
+ pkvth0 = 0 stk2 = 0 lodk2 = 1
+ steta0 = 0 lodeta0 = 1

.model phighvt_model.39 pmos
+ level = 54 lmin = 1.8E-7 lmax = 2.5E-7 wmin = 5.5E-7
+ wmax = 1E-6 version = 4.5 binunit = 2
+ mobmod = 0 capmod = 2 rdsmod = 0
+ igcmod = 0 igbmod = 0 rbodymod = 1
+ trnqsmod = 0 acnqsmod = 0 fnoimod = 1
+ tnoimod = 1 diomod = 1 tempmod = 0
+ permod = 1 geomod = 0 rgatemod = 0
+ epsrox = 3.9 toxe = 4.23E-9
+ toxm = 4.23E-9 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 9.999999999999999E22 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {9.364E-9+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {-1.176E-8-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = -5.722E-9 dwb = -1.7864E-8 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = -0.959931947413538 lvth0 = -1.783855011037123E-8
+ wvth0 = -5.807337025771501E-8 pvth0 = 9.477122194237142E-15 k1 = -2.420817069990844
+ lk1 = 7.07033393450484E-7 wk1 = 1.738566863198096E-6 pk1 = -3.756270450052255E-13
+ k2 = 1.053855865346346 lk2 = -2.507188931312642E-7 wk2 = -6.233094897422838E-7
+ pk2 = 1.33199927791633E-13 k3 = -13.778 k3b = 2
+ w0 = 0 lpe0 = 0 lpeb = 0
+ vbm = -3 dvtp0 = 0 dvtp1 = 0
+ dvt0 = 4.05 dvt1 = 0.3 dvt2 = 0.03
+ dvt0w = -4.254 dvt1w = 1.1472E6 dvt2w = -8.96E-3
+ vfbsdoff = 0 u0 = 0.031830075092685 lu0 = -5.871980846719512E-9
+ wu0 = -1.522292790912107E-8 pu0 = 2.992872406672417E-15 ua = 8.233935245517212E-9
+ lua = -2.134865841385014E-15 wua = -5.78213506893242E-15 pua = 1.134194445284299E-21
+ ub = -5.757235435363582E-18 lub = 1.563499868054281E-24 wub = 4.308650099577281E-24
+ pub = -8.30643701900934E-31 uc = 6.242499267772342E-11 luc = -1.712940154581376E-17
+ wuc = -3.302756075172748E-17 puc = 9.10037141804757E-24 ud = 0
+ up = 0 lp = 1 eu = 1.67
+ vsat = -2.752134923213596E5 lvsat = 0.10543159011028 wvsat = 0.192562985588553
+ pvsat = -5.601285174106864E-8 a0 = -2.128211188991292 la0 = 5.592310633031878E-7
+ wa0 = 1.750289517477782E-6 pa0 = -2.971038054632112E-13 ags = 3.615306375915684
+ lags = -4.813871536263603E-7 wags = -1.256621048945478E-6 pags = 2.557475158813837E-13
+ b0 = 0 b1 = 0 keta = 0.072175603354852
+ lketa = -3.049767964995243E-8 wketa = -5.333670305154702E-8 pketa = 1.620256326298953E-14
+ a1 = 0 a2 = 2.671449335949285 la2 = -3.996631871907469E-7
+ wa2 = -1.178867803260049E-6 pa2 = 2.123298607852025E-13 rdsw = 531.92
+ rdswmin = 0 rdw = 0 rdwmin = 0
+ rsw = 0 rswmin = 0 prwb = -0.32348
+ prwg = 0.02 wr = 1 voff = 0.173760249513237
+ lvoff = -9.249942596213058E-8 wvoff = -2.310917486372363E-7 pvoff = 4.914235502975304E-14
+ voffl = 0 minv = 0 nfactor = 7.254064402491594
+ lnfactor = -1.153701018852616E-6 wnfactor = -2.832478794411715E-6 pnfactor = 6.129290476878672E-13
+ eta0 = 1.01168564891415 leta0 = -1.426914586909982E-7 weta0 = -2.771569780699182E-7
+ peta0 = 7.5807976641684E-14 etab = -6.25E-6 dsub = -0.18542392186818
+ ldsub = 3.224383698327814E-7 wdsub = 4.502846901164319E-7 pdsub = -1.713024776178014E-13
+ cit = 1E-5 cdsc = 0 cdscb = 0
+ cdscd = 0 pclm = 0.130915355138428 lpclm = 7.812332578656735E-8
+ wpclm = 3.696292876999369E-7 ppclm = -4.150473553728121E-14 pdiblc1 = 0.736309991327878
+ lpdiblc1 = -1.820798353691493E-8 wpdiblc1 = -2.914249742531446E-7 ppdiblc1 = 9.673391829623868E-15
+ pdiblc2 = -8.66082676100428E-5 lpdiblc2 = 1.29158063490854E-9 wpdiblc2 = 6.981288543143124E-9
+ ppdiblc2 = -6.861806270691298E-16 pdiblcb = -0.731649142187957 lpdiblcb = 1.436559671018302E-7
+ wpdiblcb = 2.691685030684802E-7 ppdiblcb = -7.632039295412356E-14 drout = -0.115088806611822
+ ldrout = 8.700344478291883E-10 wdrout = 5.914083281358758E-7 pdrout = -4.622249411671085E-16
+ pscbe1 = 7.9996855E8 pscbe2 = 2.480047061599432E-8 lpscbe2 = -4.331885249850578E-15
+ wpscbe2 = -8.225678168614933E-15 ppscbe2 = 2.301409340458616E-21 pvag = 0
+ delta = 0.01 fprout = 0 pdits = 0
+ pditsl = 0 pditsd = 0 lambda = 0
+ vtl = 0 lc = 5E-9 xn = 3
+ alpha0 = 1E-10 alpha1 = 1E-10 beta0 = 6.905423731531409
+ lbeta0 = 5.195532127145365E-7 wbeta0 = 1.158061801145845E-6 pbeta0 = -2.760240744252772E-13
+ aigbacc = 0.43 bigbacc = 0.054 cigbacc = 0.075
+ nigbacc = 1 aigbinv = 0.35 bigbinv = 0.03
+ cigbinv = 6E-3 eigbinv = 1.1 nigbinv = 3
+ aigc = 0.43 bigc = 0.054 cigc = 0.075
+ aigsd = 0.43 bigsd = 0.054 cigsd = 0.075
+ dlcig = 0 nigc = 1 poxedge = 1
+ pigcd = 1 ntox = 1 toxref = 4.23E-9
+ agidl = -2.645202096184106E-9 lagidl = 2.161900516187012E-16 wagidl = 2.338110208608082E-15
+ pagidl = -1.148557211035706E-22 bgidl = 3.218479300986229E9 lbgidl = -451.5049073367175
+ wbgidl = -1.178615935193556E3 pbgidl = 2.398719151305926E-4 cgidl = 300
+ egidl = 0.1 noia = 1.2E41 noib = 2E25
+ noic = 0 em = 4.1E7 af = 1
+ ef = 0.88 kf = 0 lintnoi = -6E-8
+ tnoia = 1.5 tnoib = 3.5 ntnoi = 1
+ rnoia = 0.577 rnoib = 0.37 xpart = 0
+ cgso = {5.932020000000001E-11/sw_func_tox_lv_ratio} cgdo = {5.932020000000001E-11/sw_func_tox_lv_ratio} cgbo = {0/sw_func_tox_lv_ratio}
+ ckappas = 0.6 cf = 1.2E-11 clc = 1E-7
+ cle = 0.6 dlc = -2.56E-9 dwc = 0
+ vfbcv = -0.1446893 noff = 4 voffcv = -0.1375
+ acde = 0.552 moin = 14.504 cgsl = {7.513892E-12/sw_func_tox_lv_ratio}
+ cgdl = {7.513892E-12/sw_func_tox_lv_ratio} ijthsrev = 0.1 ijthsfwd = 0.1
+ xjbvs = 1 bvs = 12.8 jss = 2.17E-5
+ jsws = 8.200000000000001E-10 cjs = {7.433E-04*sw_func_psd_nw_cj} mjs = 0.34629
+ mjsws = 0.26859 cjsws = {9.2435E-11*sw_func_psd_nw_cj} cjswgs = {2.4701E-10*sw_func_psd_nw_cj}
+ mjswgs = 0.70393 pbs = 0.6587 pbsws = 0.7418
+ pbswgs = 1.3925 xrcrg1 = 12 xrcrg2 = 1
+ rbpb = 50 rbpd = 50 rbps = 50
+ rbdb = 50 rbsb = 50 gbmin = 1E-12
+ tnom = 30 ute = -5.842551717738918 lute = 1.068935226646402E-6
+ wute = 3.12656479000259E-6 pute = -5.678953557308871E-13 kt1 = -0.285596006743107
+ lkt1 = -3.637164338634162E-8 wkt1 = -1.676290629455763E-7 pkt1 = 1.932323572514849E-14
+ kt1l = 0 kt2 = -0.128821365843534 lkt2 = 1.730388089016571E-8
+ wkt2 = 4.594884709842618E-8 pkt2 = -9.193067408280119E-15 ua1 = 8.943982541608478E-10
+ lua1 = -1.661410130709865E-16 wua1 = -3.19330733524542E-16 pua1 = 8.826606829624912E-23
+ ub1 = -3.882367565169315E-18 lub1 = 9.405123883911184E-25 wub1 = 2.091586819210633E-24
+ pub1 = -4.996678976053263E-31 uc1 = -5.655969455149618E-10 luc1 = 1.187822454752328E-16
+ wuc1 = 2.578721612726248E-16 puc1 = -6.310568111811786E-23 at = 2.008582919743351E5
+ lat = -0.036193103550019 wat = -0.066843204341789 pat = 1.922838250922588E-8
+ prt = 0 njs = 1.2556 xtis = 2
+ tpb = 1.9551E-3 tpbsw = 1.4242E-4 tpbswg = 0
+ tcj = 1.2407E-3 tcjsw = 0 tcjswg = 2E-12
+ tvoff = 0 tvfbsdoff = 0 saref = 1.1E-6
+ sbref = 1.1E-6 wlod = 0 ku0 = 4.5E-8
+ kvsat = 0.4 kvth0 = 2.65E-8 tku0 = 0
+ llodku0 = 0 wlodku0 = 1 llodvth = 0
+ wlodvth = 1 lku0 = 0 wku0 = 2.5E-7
+ pku0 = 0 lkvth0 = 0 wkvth0 = 2.5E-7
+ pkvth0 = 0 stk2 = 0 lodk2 = 1
+ steta0 = 0 lodeta0 = 1

.model phighvt_model.40 pmos
+ level = 54 lmin = 1.5E-7 lmax = 1.8E-7 wmin = 5.5E-7
+ wmax = 1E-6 version = 4.5 binunit = 2
+ mobmod = 0 capmod = 2 rdsmod = 0
+ igcmod = 0 igbmod = 0 rbodymod = 1
+ trnqsmod = 0 acnqsmod = 0 fnoimod = 1
+ tnoimod = 1 diomod = 1 tempmod = 0
+ permod = 1 geomod = 0 rgatemod = 0
+ epsrox = 3.9 toxe = 4.23E-9
+ toxm = 4.23E-9 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 9.999999999999999E22 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {9.364E-9+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {-1.176E-8-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = -5.722E-9 dwb = -1.7864E-8 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = -0.468246760425753 lvth0 = -1.179063193661252E-7
+ wvth0 = -3.192919429190895E-7 pvth0 = 6.264032610228009E-14 k1 = 2.219048692624911
+ lk1 = -2.372720865570744E-7 wk1 = -7.264639002383015E-7 pk1 = 1.2605601596935E-13
+ k2 = -0.719223048905864 lk2 = 1.101381274973454E-7 wk2 = 3.18677691190316E-7
+ pk2 = -5.85133032717697E-14 k3 = -13.778 k3b = 2
+ w0 = 0 lpe0 = 0 lpeb = 0
+ vbm = -3 dvtp0 = 0 dvtp1 = 0
+ dvt0 = 4.05 dvt1 = 0.3 dvt2 = 0.03
+ dvt0w = -4.254 dvt1w = 1.1472E6 dvt2w = -8.96E-3
+ vfbsdoff = 0 u0 = 7.118912915726215E-3 lu0 = -8.427651204648125E-10
+ wu0 = -2.1027761250437E-9 pu0 = 3.226591155769902E-16 ua = 2.229926475496486E-11
+ lua = -4.636336865802814E-16 wua = -1.4195227981609E-15 pua = 2.463155959368793E-22
+ ub = -5.491852826305091E-19 lub = 5.035575009700458E-25 wub = 1.541758878834476E-24
+ pub = -2.675260006553582E-31 uc = -2.624949553054493E-10 luc = 4.899830626772155E-17
+ wuc = 1.395933098531887E-16 puc = -2.603142816746496E-23 ud = 0
+ up = 0 lp = 1 eu = 1.67
+ vsat = 1.243625421954559E6 lvsat = -0.203682505723155 wvsat = -0.614353602076642
+ pvsat = 1.08210812180552E-7 a0 = -2.542715222677329 la0 = 6.435909242389699E-7
+ wa0 = 1.97050390446223E-6 pa0 = -3.41921837502286E-13 ags = 1.25
+ b0 = 0 b1 = 0 keta = -0.666258145847802
+ lketa = 1.197883569877718E-7 wketa = 3.389724717548457E-7 pketa = -6.364019999360752E-14
+ a1 = 0 a2 = 2.183769480588384 la2 = -3.004105830276965E-7
+ wa2 = -9.197771511427525E-7 pa2 = 1.595997312662904E-13 rdsw = 531.92
+ rdswmin = 0 rdw = 0 rdwmin = 0
+ rsw = 0 rswmin = 0 prwb = -0.32348
+ prwg = 0.02 wr = 1 voff = -0.393639927559887
+ lvoff = 2.297785807579163E-8 wvoff = 7.035207823675643E-8 pvoff = -1.220749261564197E-14
+ voffl = 0 minv = 0 nfactor = -0.365217075517551
+ lnfactor = 3.969751475518052E-7 wnfactor = 1.21543211497316E-6 pnfactor = -2.109017805901427E-13
+ eta0 = -0.727266514133013 leta0 = 2.112200855323604E-7 weta0 = 6.466996154964741E-7
+ peta0 = -1.122153172809482E-13 etab = -6.25E-6 dsub = 5.660236944178967
+ ldsub = -8.672705296251343E-7 wdsub = -2.655351249510169E-6 pdsub = 4.607565488150044E-13
+ cit = 1E-5 cdsc = 0 cdscb = 0
+ cdscd = 0 pclm = -1.289156878068654 lpclm = 3.671364266888727E-7
+ wpclm = 1.12407390318033E-6 ppclm = -1.950493036798508E-13 pdiblc1 = 3.302143795404492
+ lpdiblc1 = -5.404064793425873E-7 wpdiblc1 = -1.654580631012535E-6 ppdiblc1 = 2.87102831093295E-13
+ pdiblc2 = -0.282120070438515 lpdiblc2 = 5.869103085593107E-8 wpdiblc2 = 1.56817770057604E-7
+ ppdiblc2 = -3.118090134489222E-14 pdiblcb = 1.126424456124573 lpdiblcb = -2.34499171626736E-7
+ wpdiblcb = -7.179739736542143E-7 ppdiblcb = 1.245828439084793E-13 drout = -6.524796586993618
+ ldrout = 1.305373761911132E-6 wdrout = 3.996706600034873E-6 pdrout = -6.93508529238051E-13
+ pscbe1 = 7.9996855E8 pscbe2 = -3.004209995931373E-8 lpscbe2 = 6.829674713636117E-15
+ wpscbe2 = 2.091064398607012E-14 ppscbe2 = -3.628414944462887E-21 pvag = 0
+ delta = 0.01 fprout = 0 pdits = 0
+ pditsl = 0 pditsd = 0 lambda = 0
+ vtl = 0 lc = 5E-9 xn = 3
+ alpha0 = 1E-10 alpha1 = 1E-10 beta0 = 11.615954350526955
+ lbeta0 = -4.391339788634373E-7 wbeta0 = -1.344511221869157E-6 pbeta0 = 2.332995872187361E-13
+ aigbacc = 0.43 bigbacc = 0.054 cigbacc = 0.075
+ nigbacc = 1 aigbinv = 0.35 bigbinv = 0.03
+ cigbinv = 6E-3 eigbinv = 1.1 nigbinv = 3
+ aigc = 0.43 bigc = 0.054 cigc = 0.075
+ aigsd = 0.43 bigsd = 0.054 cigsd = 0.075
+ dlcig = 0 nigc = 1 poxedge = 1
+ pigcd = 1 ntox = 1 toxref = 4.23E-9
+ agidl = -1.166706454647709E-8 lagidl = 2.052319497502329E-15 wagidl = 7.131173116300136E-15
+ pagidl = -1.090339884077058E-21 bgidl = 1E9 cgidl = 300
+ egidl = 0.1 noia = 1.2E41 noib = 2E25
+ noic = 0 em = 4.1E7 af = 1
+ ef = 0.88 kf = 0 lintnoi = -6E-8
+ tnoia = 1.5 tnoib = 3.5 ntnoi = 1
+ rnoia = 0.577 rnoib = 0.37 xpart = 0
+ cgso = {5.932020000000001E-11/sw_func_tox_lv_ratio} cgdo = {5.932020000000001E-11/sw_func_tox_lv_ratio} cgbo = {0/sw_func_tox_lv_ratio}
+ ckappas = 0.6 cf = 1.2E-11 clc = 1E-7
+ cle = 0.6 dlc = -2.56E-9 dwc = 0
+ vfbcv = -0.1446893 noff = 4 voffcv = -0.1375
+ acde = 0.552 moin = 14.504 cgsl = {7.513892E-12/sw_func_tox_lv_ratio}
+ cgdl = {7.513892E-12/sw_func_tox_lv_ratio} ijthsrev = 0.1 ijthsfwd = 0.1
+ xjbvs = 1 bvs = 12.8 jss = 2.17E-5
+ jsws = 8.200000000000001E-10 cjs = {7.433E-04*sw_func_psd_nw_cj} mjs = 0.34629
+ mjsws = 0.26859 cjsws = {9.2435E-11*sw_func_psd_nw_cj} cjswgs = {2.4701E-10*sw_func_psd_nw_cj}
+ mjswgs = 0.70393 pbs = 0.6587 pbsws = 0.7418
+ pbswgs = 1.3925 xrcrg1 = 12 xrcrg2 = 1
+ rbpb = 50 rbpd = 50 rbps = 50
+ rbdb = 50 rbsb = 50 gbmin = 1E-12
+ tnom = 30 ute = -3.020387696862575 lute = 4.945684051176482E-7
+ wute = 1.627228066303574E-6 pute = -2.627503457236632E-13 kt1 = 0.70538514057671
+ lkt1 = -2.380561264888707E-7 wkt1 = -6.941095990444698E-7 pkt1 = 1.264725544319953E-13
+ kt1l = 0 kt2 = 0.275653974562986 lkt2 = -6.501494038936934E-8
+ wkt2 = -1.689375759500268E-7 pkt2 = 3.454061741054104E-14 ua1 = -1.167056732805688E-9
+ lua1 = 2.534063058764428E-16 wua1 = 7.758625803111433E-16 pua1 = -1.346276749355895E-22
+ ub1 = 4.696775368261967E-18 lub1 = -8.055147814208164E-25 wub1 = -2.466271605319272E-24
+ pub1 = 4.27947448955E-31 uc1 = 3.104278989158573E-10 luc1 = -5.950633086332754E-17
+ wuc1 = -2.075353098778253E-16 puc1 = 3.161404741042175E-23 at = 1.323173058500976E5
+ lat = -0.022243642054015 wat = -0.030429297561593 pat = 1.181742420132041E-8
+ prt = 0 njs = 1.2556 xtis = 2
+ tpb = 1.9551E-3 tpbsw = 1.4242E-4 tpbswg = 0
+ tcj = 1.2407E-3 tcjsw = 0 tcjswg = 2E-12
+ tvoff = 0 tvfbsdoff = 0 saref = 1.1E-6
+ sbref = 1.1E-6 wlod = 0 ku0 = 4.5E-8
+ kvsat = 0.4 kvth0 = 2.65E-8 tku0 = 0
+ llodku0 = 0 wlodku0 = 1 llodvth = 0
+ wlodvth = 1 lku0 = 0 wku0 = 2.5E-7
+ pku0 = 0 lkvth0 = 0 wkvth0 = 2.5E-7
+ pkvth0 = 0 stk2 = 0 lodk2 = 1
+ steta0 = 0 lodeta0 = 1

.model phighvt_model.41 pmos
+ level = 54 lmin = 8E-6 lmax = 2.02E-5 wmin = 4.2E-7
+ wmax = 5.5E-7 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 4.23E-9
+ toxm = 4.23E-9 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 9.999999999999999E22 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {9.364E-9+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {-1.176E-8-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = -5.722E-9 dwb = -1.7864E-8 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = -0.874646958222745 lvth0 = -1.037686905196761E-6
+ wvth0 = -1.077231767662859E-7 pvth0 = 5.512939974976936E-13 k1 = 0.520628336754318
+ lk1 = 6.93609598439888E-9 wk1 = -3.565723234350022E-8 pk1 = -3.684953585823562E-15
+ k2 = 0.029400031717085 lk2 = -2.033313810333703E-7 wk2 = -2.291182071415106E-9
+ pk2 = 1.080242694643607E-13 k3 = -13.778 k3b = 2
+ w0 = 0 lpe0 = 0 lpeb = 0
+ vbm = -3 dvtp0 = 0 dvtp1 = 0
+ dvt0 = 4.05 dvt1 = 0.3 dvt2 = 0.03
+ dvt0w = -4.254 dvt1w = 1.1472E6 dvt2w = -8.96E-3
+ vfbsdoff = 0 u0 = 1.423140747667437E-3 lu0 = 4.400519809357705E-8
+ wu0 = 3.561385173689226E-9 pu0 = -2.337872960157086E-14 ua = 6.346357780223614E-10
+ lua = -7.59787946510346E-15 wua = -6.039723591623761E-16 pua = 4.036540619184446E-21
+ ub = -2.461438695039239E-18 lub = 2.068870228592711E-23 wub = 1.503419604357847E-24
+ pub = -1.099132824084907E-29 uc = -1.205936282360252E-10 luc = 1.754141319295339E-16
+ wuc = 7.130099633169561E-18 puc = -9.319261669846734E-23 ud = 0
+ up = 0 lp = 1 eu = 1.67
+ vsat = 2.132593085292334E3 wvsat = 0.031308608539479 a0 = 0.330676580745108
+ la0 = 2.801878620961383E-6 wa0 = 4.729617737247848E-7 pa0 = -1.488559658715396E-12
+ ags = 0.142179488617838 lags = -5.116114650074042E-7 wags = -1.4914111234816E-8
+ pags = 2.718048462374137E-13 b0 = 4.907812258307558E-7 lb0 = -2.572851905365991E-12
+ wb0 = -2.488001102975573E-13 pb0 = 1.366884177467601E-18 b1 = 3.494401684152914E-8
+ lb1 = -2.792762927894E-13 wb1 = -1.854926244794488E-14 pb1 = 1.483716746228102E-19
+ keta = -0.04086014214278 lketa = -4.224232879840051E-8 wketa = 2.549599746325238E-8
+ pketa = 2.244216650538384E-14 a1 = 0 a2 = 0.275259692307693
+ wa2 = 2.787798327483075E-7 rdsw = 531.92 rdswmin = 0
+ rdw = 0 rdwmin = 0 rsw = 0
+ rswmin = 0 prwb = -0.32348 prwg = 0.02
+ wr = 1 voff = -0.04266247379509 lvoff = -1.544225647479639E-6
+ wvoff = -8.540672686817504E-8 pvoff = 8.204038481878028E-13 voffl = 0
+ minv = 0 nfactor = 1.953882328251692 lnfactor = -3.339085949707213E-5
+ wnfactor = -2.476800308261328E-7 pnfactor = 1.773962870672851E-11 eta0 = 0.08
+ etab = -0.07 dsub = 0.56 cit = 5.983346049235874E-5
+ lcit = -3.998397669296502E-10 wcit = -2.647512222269641E-11 pcit = 2.124236726562491E-16
+ cdsc = 0 cdscb = 0 cdscd = 0
+ pclm = 0.534715622338204 lpclm = -9.92784114129037E-8 wpclm = -2.091918788883023E-7
+ ppclm = 5.274384018815617E-14 pdiblc1 = 0.39 pdiblc2 = 1.146002990131838E-3
+ lpdiblc2 = -7.477997906231086E-8 wpdiblc2 = -4.328697630410014E-10 ppdiblc2 = 3.972850903639201E-14
+ pdiblcb = -0.225 drout = 0.56 pscbe1 = 5.111619962386229E8
+ lpscbe1 = 5.78355354507601E3 wpscbe1 = 153.45154393431434 ppscbe1 = -3.072640058999622E-3
+ pscbe2 = 1.666711338806459E-8 lpscbe2 = 1.455976389073762E-14 wpscbe2 = -2.556471507271853E-15
+ ppscbe2 = -7.735194881759955E-21 pvag = 0 delta = 0.01
+ fprout = 0 pdits = 0 pditsl = 0
+ pditsd = 0 lambda = 0 vtl = 0
+ lc = 5E-9 xn = 3 alpha0 = 4.086707692307691E-10
+ walpha0 = -1.639881369107692E-16 alpha1 = 4.086707692307691E-10 walpha1 = -1.639881369107692E-16
+ beta0 = -80.34110769230766 wbeta0 = 4.427679696590768E-5 aigbacc = 0.43
+ bigbacc = 0.054 cigbacc = 0.075 nigbacc = 1
+ aigbinv = 0.35 bigbinv = 0.03 cigbinv = 6E-3
+ eigbinv = 1.1 nigbinv = 3 aigc = 0.43
+ bigc = 0.054 cigc = 0.075 aigsd = 0.43
+ bigsd = 0.054 cigsd = 0.075 dlcig = 0
+ nigc = 1 poxedge = 1 pigcd = 1
+ ntox = 1 toxref = 4.23E-9 agidl = -6.045779404465611E-9
+ lagidl = 4.752959608005905E-14 wagidl = 3.497101565647494E-15 pagidl = -2.525114356864513E-20
+ bgidl = 1E9 cgidl = 300 egidl = 0.1
+ noia = 1.2E41 noib = 2E25 noic = 0
+ em = 4.1E7 af = 1 ef = 0.88
+ kf = 0 lintnoi = -6E-8 tnoia = 1.5
+ tnoib = 3.5 ntnoi = 1 rnoia = 0.577
+ rnoib = 0.37 xpart = 0 cgso = {5.932020000000001E-11/sw_func_tox_lv_ratio}
+ cgdo = {5.932020000000001E-11/sw_func_tox_lv_ratio} cgbo = {0/sw_func_tox_lv_ratio} ckappas = 0.6
+ cf = 1.2E-11 clc = 1E-7 cle = 0.6
+ dlc = -2.56E-9 dwc = 0 vfbcv = -0.1446893
+ noff = 4 voffcv = -0.1375 acde = 0.552
+ moin = 14.504 cgsl = {7.513892E-12/sw_func_tox_lv_ratio} cgdl = {7.513892E-12/sw_func_tox_lv_ratio}
+ ijthsrev = 0.1 ijthsfwd = 0.1 xjbvs = 1
+ bvs = 12.8 jss = 2.17E-5 jsws = 8.200000000000001E-10
+ cjs = {7.433E-04*sw_func_psd_nw_cj} mjs = 0.34629 mjsws = 0.26859
+ cjsws = {9.2435E-11*sw_func_psd_nw_cj} cjswgs = {2.4701E-10*sw_func_psd_nw_cj} mjswgs = 0.70393
+ pbs = 0.6587 pbsws = 0.7418 pbswgs = 1.3925
+ xrcrg1 = 12 xrcrg2 = 1 rbpb = 50
+ rbpd = 50 rbps = 50 rbdb = 50
+ rbsb = 50 gbmin = 1E-12 tnom = 30
+ ute = -5.99407649145777 lute = 3.938003208682193E-5 wute = 2.627627052504153E-6
+ pute = -2.092150840683006E-11 kt1 = -0.540621262855524 lkt1 = 2.801465364527622E-6
+ wkt1 = 5.926685701050009E-8 pkt1 = -1.488340107143319E-12 kt1l = 0
+ kt2 = -4.697481315533963E-3 lkt2 = -2.610127635692056E-7 wkt2 = -2.330249291476564E-8
+ pkt2 = 1.38668772926939E-13 ua1 = -1.152226846058602E-8 lua1 = 6.630782131128273E-14
+ wua1 = 5.892797021017173E-15 pua1 = -3.52274888436878E-20 ub1 = 9.424942810171515E-18
+ lub1 = -3.953748278808836E-23 wub1 = -4.531780580725842E-24 pub1 = 2.100515755579328E-29
+ uc1 = 5.345211467783489E-10 luc1 = -3.385851287521941E-15 wuc1 = -2.48424043540523E-16
+ puc1 = 1.798807985224356E-21 at = -9.259770990994453E4 lat = 2.52045098956394
+ wat = 0.082006855266372 pat = -1.339045038127614E-6 prt = 0
+ njs = 1.2556 xtis = 2 tpb = 1.9551E-3
+ tpbsw = 1.4242E-4 tpbswg = 0 tcj = 1.2407E-3
+ tcjsw = 0 tcjswg = 2E-12 tvoff = 0
+ tvfbsdoff = 0 saref = 3E-6 sbref = 3E-6
+ wlod = 0 ku0 = 4.5E-8 kvsat = 0.4
+ kvth0 = 2.65E-8 tku0 = 0 llodku0 = 0
+ wlodku0 = 1 llodvth = 0 wlodvth = 1
+ lku0 = 0 wku0 = 2.5E-7 pku0 = 0
+ lkvth0 = 0 wkvth0 = 2.5E-7 pkvth0 = 0
+ stk2 = 0 lodk2 = 1 steta0 = 0
+ lodeta0 = 1

.model phighvt_model.42 pmos
+ level = 54 lmin = 4E-6 lmax = 8E-6 wmin = 4.2E-7
+ wmax = 5.5E-7 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 4.23E-9
+ toxm = 4.23E-9 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 9.999999999999999E22 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {9.364E-9+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {-1.176E-8-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = -5.722E-9 dwb = -1.7864E-8 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = -0.965942647972967 lvth0 = -3.051741125720624E-7
+ wvth0 = -4.49870194720801E-8 pvth0 = 4.792918472448765E-14 k1 = 0.519617777016782
+ lk1 = 1.504434224971255E-8 wk1 = -3.145526023953504E-8 pk1 = -3.739956080143029E-14
+ k2 = 0.019247760150652 lk2 = -1.218744270746666E-7 wk2 = 6.304078748874962E-9
+ pk2 = 3.906002236754691E-14 k3 = -13.778 k3b = 2
+ w0 = 0 lpe0 = 0 lpeb = 0
+ vbm = -3 dvtp0 = 0 dvtp1 = 0
+ dvt0 = 4.05 dvt1 = 0.3 dvt2 = 0.03
+ dvt0w = -4.254 dvt1w = 1.1472E6 dvt2w = -8.96E-3
+ vfbsdoff = 0 u0 = 3.093826836193176E-3 lu0 = 3.060041484856901E-8
+ wu0 = 1.331144956633878E-9 pu0 = -5.484352615222941E-15 ua = -4.704338238773036E-10
+ lua = 1.26866858713054E-15 wua = -2.798077912825328E-17 pua = -5.84939343050939E-22
+ ub = -4.424126262097877E-19 lub = 4.489006242152624E-24 wub = 1.931199810048513E-25
+ pub = -4.781130068838387E-31 uc = -8.938960222025083E-11 luc = -7.495199488855188E-17
+ wuc = -9.359683955158351E-18 puc = 3.911349171815344E-23 ud = 0
+ up = 0 lp = 1 eu = 1.67
+ vsat = -6.684254095868117E4 lvsat = 0.553423367504502 wvsat = 0.069216004871742
+ pvsat = -3.041507526198445E-7 a0 = 0.043892649186151 la0 = 5.102895231503313E-6
+ wa0 = 5.978458152767413E-7 pa0 = -2.490569263788351E-12 ags = 4.367968379367204E-3
+ lags = 5.941220238563704E-7 wags = 2.146333604481408E-8 pags = -2.007032955964385E-14
+ b0 = 4.690374859087629E-7 lb0 = -2.398390573227082E-12 wb0 = -1.878781067870467E-13
+ pb0 = 8.780752638609484E-19 b1 = -7.316223698170802E-9 lb1 = 5.979959238569336E-14
+ wb1 = 3.809260967997288E-15 pb1 = -3.102238517547014E-20 keta = -0.07779191854544
+ lketa = 2.540805178038744E-7 wketa = 4.53346717946373E-8 pketa = -1.367338337659696E-13
+ a1 = 0 a2 = -0.252566088393845 la2 = 4.235020707974405E-6
+ wa2 = 5.59198890913175E-7 pa2 = -2.249947921566978E-12 rdsw = 531.92
+ rdswmin = 0 rdw = 0 rdwmin = 0
+ rsw = 0 rswmin = 0 prwb = -0.32348
+ prwg = 0.02 wr = 1 voff = -0.285954688637776
+ lvoff = 4.078343041549516E-7 wvoff = 5.08086340444368E-8 pvoff = -2.725228244017566E-13
+ voffl = 0 minv = 0 nfactor = -7.4502731705679
+ lnfactor = 4.206357023081684E-5 wnfactor = 4.371559237512113E-6 pnfactor = -1.932292994756878E-11
+ eta0 = 0.08 etab = -0.07 dsub = 0.56
+ cit = 1E-5 cdsc = 0 cdscb = 0
+ cdscd = 0 pclm = -0.72199746722876 lpclm = 9.983984196989422E-6
+ wpclm = 1.652595022650794E-7 ppclm = -2.951674305523625E-12 pdiblc1 = 0.39
+ pdiblc2 = -0.016367560887872 lpdiblc2 = 6.574045098412846E-8 wpdiblc2 = 8.81881035584193E-9
+ ppdiblc2 = -3.450253143106755E-14 pdiblcb = -0.225 drout = 0.56
+ pscbe1 = 1.666514011284132E9 lpscbe1 = -3.486436454681929E3 wpscbe1 = -460.3546318029432
+ ppscbe1 = 1.852246068151778E-3 pscbe2 = 2.935529764311571E-8 lpscbe2 = -8.724413624335015E-14
+ wpscbe2 = -7.820535633886244E-15 ppscbe2 = 3.450112891941315E-20 pvag = 0
+ delta = 0.01 fprout = 0 pdits = 0
+ pditsl = 0 pditsd = 0 lambda = 0
+ vtl = 0 lc = 5E-9 xn = 3
+ alpha0 = 8.197445225846151E-10 lalpha0 = -3.298258481509651E-15 walpha0 = -3.289405240665737E-16
+ palpha0 = 1.32349877739234E-21 alpha1 = 8.197445225846151E-10 lalpha1 = -3.298258481509651E-15
+ walpha1 = -3.289405240665737E-16 palpha1 = 1.32349877739234E-21 beta0 = -191.3310210978461
+ lbeta0 = 8.905297900076057E-4 wbeta0 = 8.88139414979749E-5 pbeta0 = -3.573446698959319E-10
+ aigbacc = 0.43 bigbacc = 0.054 cigbacc = 0.075
+ nigbacc = 1 aigbinv = 0.35 bigbinv = 0.03
+ cigbinv = 6E-3 eigbinv = 1.1 nigbinv = 3
+ aigc = 0.43 bigc = 0.054 cigc = 0.075
+ aigsd = 0.43 bigsd = 0.054 cigsd = 0.075
+ dlcig = 0 nigc = 1 poxedge = 1
+ pigcd = 1 ntox = 1 toxref = 4.23E-9
+ agidl = 2.77102634172688E-9 lagidl = -2.321222116063133E-14 wagidl = -1.10312877920281E-15
+ pagidl = 1.165889660786818E-20 bgidl = 1E9 cgidl = 300
+ egidl = 0.1 noia = 1.2E41 noib = 2E25
+ noic = 0 em = 4.1E7 af = 1
+ ef = 0.88 kf = 0 lintnoi = -6E-8
+ tnoia = 1.5 tnoib = 3.5 ntnoi = 1
+ rnoia = 0.577 rnoib = 0.37 xpart = 0
+ cgso = {5.932020000000001E-11/sw_func_tox_lv_ratio} cgdo = {5.932020000000001E-11/sw_func_tox_lv_ratio} cgbo = {0/sw_func_tox_lv_ratio}
+ ckappas = 0.6 cf = 1.2E-11 clc = 1E-7
+ cle = 0.6 dlc = -2.56E-9 dwc = 0
+ vfbcv = -0.1446893 noff = 4 voffcv = -0.1375
+ acde = 0.552 moin = 14.504 cgsl = {7.513892E-12/sw_func_tox_lv_ratio}
+ cgdl = {7.513892E-12/sw_func_tox_lv_ratio} ijthsrev = 0.1 ijthsfwd = 0.1
+ xjbvs = 1 bvs = 12.8 jss = 2.17E-5
+ jsws = 8.200000000000001E-10 cjs = {7.433E-04*sw_func_psd_nw_cj} mjs = 0.34629
+ mjsws = 0.26859 cjsws = {9.2435E-11*sw_func_psd_nw_cj} cjswgs = {2.4701E-10*sw_func_psd_nw_cj}
+ mjswgs = 0.70393 pbs = 0.6587 pbsws = 0.7418
+ pbswgs = 1.3925 xrcrg1 = 12 xrcrg2 = 1
+ rbpb = 50 rbpd = 50 rbps = 50
+ rbdb = 50 rbsb = 50 gbmin = 1E-12
+ tnom = 30 ute = -1.808042756567521 lute = 5.793306694255321E-6
+ wute = -5.864398192396885E-8 pute = 6.318409633246583E-13 kt1 = 0.143533448267266
+ lkt1 = -2.687863643260311E-6 wkt1 = -2.960904443061169E-7 pkt1 = 1.362876307116584E-12
+ kt1l = 0 kt2 = -0.015785524233505 lkt2 = -1.720476294560093E-7
+ wkt2 = -1.207481125613536E-8 pkt2 = 4.858324458528572E-14 ua1 = -8.637822907899594E-9
+ lua1 = 4.316441473039218E-14 wua1 = 3.013371477595978E-15 pua1 = -1.212436040753697E-20
+ ub1 = 1.015647151904475E-17 lub1 = -4.540691801430695E-23 wub1 = -3.838918642318034E-24
+ pub1 = 1.544596593573945E-29 uc1 = 1.852095647226464E-9 luc1 = -1.39574366433574E-14
+ wuc1 = -6.892010691944134E-16 puc1 = 5.33539126609886E-21 at = 2.496433058306716E5
+ lat = -0.225526645051209 wat = -0.120779632543452 pat = 2.880164025442633E-7
+ prt = 0 njs = 1.2556 xtis = 2
+ tpb = 1.9551E-3 tpbsw = 1.4242E-4 tpbswg = 0
+ tcj = 1.2407E-3 tcjsw = 0 tcjswg = 2E-12
+ tvoff = 0 tvfbsdoff = 0 saref = 3E-6
+ sbref = 3E-6 wlod = 0 ku0 = 4.5E-8
+ kvsat = 0.4 kvth0 = 2.65E-8 tku0 = 0
+ llodku0 = 0 wlodku0 = 1 llodvth = 0
+ wlodvth = 1 lku0 = 0 wku0 = 2.5E-7
+ pku0 = 0 lkvth0 = 0 wkvth0 = 2.5E-7
+ pkvth0 = 0 stk2 = 0 lodk2 = 1
+ steta0 = 0 lodeta0 = 1

.model phighvt_model.43 pmos
+ level = 54 lmin = 2E-6 lmax = 4E-6 wmin = 4.2E-7
+ wmax = 5.5E-7 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 4.23E-9
+ toxm = 4.23E-9 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 9.999999999999999E22 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {9.364E-9+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {-1.176E-8-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = -5.722E-9 dwb = -1.7864E-8 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = -0.917053016403955 lvth0 = -5.0188252298261E-7
+ wvth0 = -1.004500295326283E-7 pvth0 = 2.710857149633047E-13 k1 = 0.42904626660568
+ lk1 = 3.794606258189908E-7 wk1 = -2.321926139663938E-8 pk1 = -7.053726686579784E-14
+ k2 = 0.067628109875306 lk2 = -3.16533731798806E-7 wk2 = -1.433298360537502E-8
+ pk2 = 1.220936554911188E-13 k3 = -13.778 k3b = 2
+ w0 = 0 lpe0 = 0 lpeb = 0
+ vbm = -3 dvtp0 = 0 dvtp1 = 0
+ dvt0 = 4.05 dvt1 = 0.3 dvt2 = 0.03
+ dvt0w = -4.254 dvt1w = 1.1472E6 dvt2w = -8.96E-3
+ vfbsdoff = 0 u0 = 3.160011138617153E-3 lu0 = 3.033412098408008E-8
+ wu0 = 4.75682568821598E-9 pu0 = -1.926764755235816E-14 ua = -2.067684362209853E-10
+ lua = 2.078056265875907E-16 wua = 4.032625991665658E-17 pua = -8.597740807889148E-22
+ ub = -5.84896664505419E-19 lub = 5.062293619915861E-24 wub = 6.39463023729089E-25
+ pub = -2.273983166145663E-30 uc = -9.733710513792727E-11 luc = -4.297505794922229E-17
+ wuc = -1.937642430264727E-17 puc = 7.941604684108207E-23 ud = 0
+ up = 0 lp = 1 eu = 1.67
+ vsat = 1.608224484151262E5 lvsat = -0.362591270540799 wvsat = -0.040872292865193
+ pvsat = 1.387917150906694E-7 a0 = 1.744050646939864 la0 = -1.737724475618711E-6
+ wa0 = -1.823779620578021E-7 pa0 = 6.486767087927316E-13 ags = -0.506336178152166
+ lags = 2.648950371508922E-6 wags = 2.454557399006112E-7 pags = -9.213082463215208E-13
+ b0 = -2.77108107760936E-8 lb0 = -3.997138665496278E-13 wb0 = -3.861738059535553E-14
+ pb0 = 2.77521746814155E-19 b1 = 2.168399396965884E-8 lb1 = -5.68833634051725E-14
+ wb1 = -1.04623167707652E-14 pb1 = 2.63995932879955E-20 keta = 5.144175734482452E-3
+ lketa = -7.96145162532796E-8 wketa = 9.385855764138204E-9 pketa = 7.906946509064061E-15
+ a1 = 0 a2 = 0.8 rdsw = 531.92
+ rdswmin = 0 rdw = 0 rdwmin = 0
+ rsw = 0 rswmin = 0 prwb = -0.32348
+ prwg = 0.02 wr = 1 voff = -0.033714237461816
+ lvoff = -6.070601959605491E-7 wvoff = -1.002285081769047E-7 pvoff = 3.351781380686555E-13
+ voffl = 0 minv = 0 nfactor = 6.391607816008558
+ lnfactor = -1.362951475629327E-5 wnfactor = -2.189183389064302E-6 pnfactor = 7.074349225313964E-12
+ eta0 = 0.16043492 leta0 = -3.236315093184E-7 etab = -0.14031732
+ letab = 2.829231433664E-7 dsub = 0.863527958652327 ldsub = -1.221250812196809E-6
+ pdsub = -6.675689048578964E-20 cit = 1E-5 cdsc = 0
+ cdscb = 0 cdscd = 0 pclm = 2.32889232220562
+ lpclm = -2.291331888595596E-6 wpclm = -9.153296284845989E-7 ppclm = 1.39609767383032E-12
+ pdiblc1 = 0.39 pdiblc2 = -5.3925634099929E-4 lpdiblc2 = 2.054951073696189E-9
+ wpdiblc2 = 5.088520584291498E-10 ppdiblc2 = -1.067248022261289E-15 pdiblcb = -1.051953474953846
+ lpdiblcb = 3.327263845546298E-6 wpdiblcb = 3.318332748016797E-7 ppdiblcb = -1.335137817830054E-12
+ drout = 0.56 pscbe1 = 8E8 pscbe2 = 5.580637980926026E-9
+ lpscbe2 = 8.413682400663303E-15 wpscbe2 = 1.663859180567648E-15 ppscbe2 = -3.659523304438379E-21
+ pvag = 0 delta = 0.01 fprout = 0
+ pdits = 0 pditsl = 0 pditsd = 0
+ lambda = 0 vtl = 0 lc = 5E-9
+ xn = 3 alpha0 = -1.01176E-10 lalpha0 = 4.0708365952E-16
+ alpha1 = -1.01176E-10 lalpha1 = 4.0708365952E-16 beta0 = 51.75207830848191
+ lbeta0 = -8.751992211574316E-5 wbeta0 = 1.576468876261972E-6 pbeta0 = -6.342954053017569E-12
+ aigbacc = 0.43 bigbacc = 0.054 cigbacc = 0.075
+ nigbacc = 1 aigbinv = 0.35 bigbinv = 0.03
+ cigbinv = 6E-3 eigbinv = 1.1 nigbinv = 3
+ aigc = 0.43 bigc = 0.054 cigc = 0.075
+ aigsd = 0.43 bigsd = 0.054 cigsd = 0.075
+ dlcig = 0 nigc = 1 poxedge = 1
+ pigcd = 1 ntox = 1 toxref = 4.23E-9
+ agidl = -3.336956655430773E-9 lagidl = 1.363370588092429E-15 wagidl = 1.733787257832962E-15
+ pagidl = 2.445081945340147E-22 bgidl = 1E9 cgidl = 300
+ egidl = 0.1 noia = 1.2E41 noib = 2E25
+ noic = 0 em = 4.1E7 af = 1
+ ef = 0.88 kf = 0 lintnoi = -6E-8
+ tnoia = 1.5 tnoib = 3.5 ntnoi = 1
+ rnoia = 0.577 rnoib = 0.37 xpart = 0
+ cgso = {5.932020000000001E-11/sw_func_tox_lv_ratio} cgdo = {5.932020000000001E-11/sw_func_tox_lv_ratio} cgbo = {0/sw_func_tox_lv_ratio}
+ ckappas = 0.6 cf = 1.2E-11 clc = 1E-7
+ cle = 0.6 dlc = -2.56E-9 dwc = 0
+ vfbcv = -0.1446893 noff = 4 voffcv = -0.1375
+ acde = 0.552 moin = 14.504 cgsl = {7.513892E-12/sw_func_tox_lv_ratio}
+ cgdl = {7.513892E-12/sw_func_tox_lv_ratio} ijthsrev = 0.1 ijthsfwd = 0.1
+ xjbvs = 1 bvs = 12.8 jss = 2.17E-5
+ jsws = 8.200000000000001E-10 cjs = {7.433E-04*sw_func_psd_nw_cj} mjs = 0.34629
+ mjsws = 0.26859 cjsws = {9.2435E-11*sw_func_psd_nw_cj} cjswgs = {2.4701E-10*sw_func_psd_nw_cj}
+ mjswgs = 0.70393 pbs = 0.6587 pbsws = 0.7418
+ pbswgs = 1.3925 xrcrg1 = 12 xrcrg2 = 1
+ rbpb = 50 rbpd = 50 rbps = 50
+ rbdb = 50 rbsb = 50 gbmin = 1E-12
+ tnom = 30 ute = -2.939269647697969 lute = 1.03448207152565E-5
+ wute = 1.512915174307322E-6 pute = -5.691358732955064E-12 kt1 = -0.856721743903557
+ lkt1 = 1.336683127542839E-6 wkt1 = 2.237681086472968E-7 pkt1 = -7.287849778625349E-13
+ kt1l = 0 kt2 = -0.057886497786018 lkt2 = -2.653520347998949E-9
+ wkt2 = -2.828878667684316E-9 pkt2 = 1.13820498970012E-14 ua1 = 2.417112934229674E-10
+ lua1 = 7.437431280686823E-15 wua1 = 1.405347102112594E-15 pua1 = -5.654442172292062E-21
+ ub1 = -1.62427899152448E-18 lub1 = 1.993167279978578E-24 wub1 = -1.490429153771742E-25
+ pub1 = 5.99677150878368E-31 uc1 = -3.236798277635224E-9 luc1 = 6.517829841202096E-15
+ wuc1 = 1.253619781616353E-15 puc1 = -2.481587283555276E-21 at = 2.551248129394904E5
+ lat = -0.247581598533683 wat = -0.049126756085522 pat = -2.803789417443113E-10
+ prt = 0 njs = 1.2556 xtis = 2
+ tpb = 1.9551E-3 tpbsw = 1.4242E-4 tpbswg = 0
+ tcj = 1.2407E-3 tcjsw = 0 tcjswg = 2E-12
+ tvoff = 0 tvfbsdoff = 0 saref = 3E-6
+ sbref = 3E-6 wlod = 0 ku0 = 4.5E-8
+ kvsat = 0.4 kvth0 = 2.65E-8 tku0 = 0
+ llodku0 = 0 wlodku0 = 1 llodvth = 0
+ wlodvth = 1 lku0 = 0 wku0 = 2.5E-7
+ pku0 = 0 lkvth0 = 0 wkvth0 = 2.5E-7
+ pkvth0 = 0 stk2 = 0 lodk2 = 1
+ steta0 = 0 lodeta0 = 1

.model phighvt_model.44 pmos
+ level = 54 lmin = 1E-6 lmax = 2E-6 wmin = 4.2E-7
+ wmax = 5.5E-7 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 4.23E-9
+ toxm = 4.23E-9 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 9.999999999999999E22 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {9.364E-9+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {-1.176E-8-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = -5.722E-9 dwb = -1.7864E-8 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = -1.329104455971975 lvth0 = 3.319118060120693E-7
+ wvth0 = 1.12097261676305E-7 pvth0 = -1.590079797437961E-13 k1 = 0.641442402530837
+ lk1 = -5.032720314828279E-8 wk1 = -7.170958337062879E-8 pk1 = 2.758386945500924E-14
+ k2 = -0.143682539421556 lk2 = 1.110575932663809E-7 wk2 = 7.486836336840682E-8
+ pk2 = -5.840705413726817E-14 k3 = -13.778 k3b = 2
+ w0 = 0 lpe0 = 0 lpeb = 0
+ vbm = -3 dvtp0 = 0 dvtp1 = 0
+ dvt0 = 4.05 dvt1 = 0.3 dvt2 = 0.03
+ dvt0w = -4.254 dvt1w = 1.1472E6 dvt2w = -8.96E-3
+ vfbsdoff = 0 u0 = 0.031964335301179 lu0 = -2.795200504534743E-8
+ wu0 = -1.089385515981409E-8 pu0 = 1.240181815724765E-14 ua = 1.36238396861836E-9
+ lua = -2.96740564765292E-15 wua = -9.000932778092508E-16 pua = 1.043183662190213E-21
+ ub = 2.438105245992518E-18 lub = -1.054811206014925E-24 wub = -9.164751599219774E-25
+ pub = 8.744888672359424E-31 uc = -2.281603108205428E-10 luc = 2.21748315213664E-16
+ wuc = 5.765010266785331E-17 puc = -7.644867101426528E-23 ud = 0
+ up = 0 lp = 1 eu = 1.67
+ vsat = -1.267150323942878E5 lvsat = 0.219246572626666 wvsat = 0.075487896923364
+ pvsat = -9.66654561502725E-8 a0 = 0.101369460770212 la0 = 1.586273758219305E-6
+ wa0 = 4.938540186413519E-7 pa0 = -7.196922287916204E-13 ags = 1.801743026310874
+ lags = -2.021494060306128E-6 wags = -8.256893023869184E-7 pags = 1.246175169648141E-12
+ b0 = -2.657324573080811E-7 lb0 = 8.192769564077952E-14 wb0 = 1.494279917955062E-13
+ pb0 = -1.029918251262016E-19 b1 = -1.19190227867718E-8 lb1 = 1.111301306179999E-14
+ wb1 = 4.719559985086735E-15 pb1 = -4.321237965006007E-21 keta = -0.108732006344483
+ lketa = 1.508162157071485E-7 wketa = 4.846272882254914E-8 pketa = -7.116588766209163E-14
+ a1 = 0 a2 = 0.8 rdsw = 531.92
+ rdswmin = 0 rdw = 0 rdwmin = 0
+ rsw = 0 rswmin = 0 prwb = -0.32348
+ prwg = 0.02 wr = 1 voff = -0.425236773979849
+ lvoff = 1.851934871344208E-7 wvoff = 1.168773980634238E-7 pvoff = -1.041400053267742E-13
+ voffl = 0 minv = 0 nfactor = 0.652801271453892
+ lnfactor = -2.016924937256012E-6 wnfactor = 9.856835522271465E-7 pnfactor = 6.499424722718916E-13
+ eta0 = -1.353525945452307 leta0 = 2.739898581141652E-6 weta0 = 4.531818723054581E-7
+ peta0 = -9.170225822475408E-13 etab = -2.669724509860045 letab = 5.401229180191997E-6
+ wetab = 1.418490423619301E-6 petab = -2.870343742002128E-12 dsub = 2.597887305046114
+ ldsub = -4.730761636811566E-6 wdsub = -1.242054053576064E-6 pdsub = 2.513321185308911E-12
+ cit = 1E-5 cdsc = 0 cdscb = 0
+ cdscd = 0 pclm = 1.064008530181907 lpclm = 2.681857622402289E-7
+ wpclm = -7.655157678354809E-8 ppclm = -3.011864893477898E-13 pdiblc1 = 0.40941146985677
+ lpdiblc1 = -3.927949748457101E-8 wpdiblc1 = -7.23457862497046E-9 ppdiblc1 = 1.463931453920023E-14
+ pdiblc2 = 5.236414825573063E-4 lpdiblc2 = -9.584393022705415E-11 wpdiblc2 = -3.757570498873542E-11
+ ppdiblc2 = 3.845948557007048E-17 pdiblcb = 1.428906949907692 lpdiblcb = -1.69280684136952E-6
+ wpdiblcb = -6.636665496033592E-7 ppdiblcb = 6.792759868500302E-13 drout = 0.721946231938161
+ ldrout = -3.27701439251508E-7 wdrout = -1.819393123182895E-7 pdrout = 3.681578372623053E-13
+ pscbe1 = 8E8 pscbe2 = 1.008442910008288E-8 lpscbe2 = -6.998290047729732E-16
+ wpscbe2 = -1.67299049628515E-16 ppscbe2 = 4.586199752816029E-23 pvag = 0
+ delta = 0.01 fprout = 0 pdits = 0
+ pditsl = 0 pditsd = 0 lambda = 0
+ vtl = 0 lc = 5E-9 xn = 3
+ alpha0 = 2.700078259452599E-11 lalpha0 = 1.477153764043248E-16 walpha0 = 3.878244022944099E-17
+ palpha0 = -7.847704345307842E-23 alpha1 = -5.318614114461533E-10 lalpha1 = 1.27858420328952E-15
+ walpha1 = 3.356902757818208E-16 palpha1 = -6.792759868500302E-22 beta0 = 9.912712964206946
+ lbeta0 = -2.857129554295879E-6 wbeta0 = -2.799522862335705E-6 pbeta0 = 2.511952749869603E-12
+ aigbacc = 0.43 bigbacc = 0.054 cigbacc = 0.075
+ nigbacc = 1 aigbinv = 0.35 bigbinv = 0.03
+ cigbinv = 6E-3 eigbinv = 1.1 nigbinv = 3
+ aigc = 0.43 bigc = 0.054 cigc = 0.075
+ aigsd = 0.43 bigsd = 0.054 cigsd = 0.075
+ dlcig = 0 nigc = 1 poxedge = 1
+ pigcd = 1 ntox = 1 toxref = 4.23E-9
+ agidl = -7.095585819813296E-9 lagidl = 8.969031874803749E-15 wagidl = 3.988441101171508E-15
+ pagidl = -4.3178289505384E-21 bgidl = 1E9 cgidl = 300
+ egidl = 0.1 noia = 1.2E41 noib = 2E25
+ noic = 0 em = 4.1E7 af = 1
+ ef = 0.88 kf = 0 lintnoi = -6E-8
+ tnoia = 1.5 tnoib = 3.5 ntnoi = 1
+ rnoia = 0.577 rnoib = 0.37 xpart = 0
+ cgso = {5.932020000000001E-11/sw_func_tox_lv_ratio} cgdo = {5.932020000000001E-11/sw_func_tox_lv_ratio} cgbo = {0/sw_func_tox_lv_ratio}
+ ckappas = 0.6 cf = 1.2E-11 clc = 1E-7
+ cle = 0.6 dlc = -2.56E-9 dwc = 0
+ vfbcv = -0.1446893 noff = 4 voffcv = -0.1375
+ acde = 0.552 moin = 14.504 cgsl = {7.513892E-12/sw_func_tox_lv_ratio}
+ cgdl = {7.513892E-12/sw_func_tox_lv_ratio} ijthsrev = 0.1 ijthsfwd = 0.1
+ xjbvs = 1 bvs = 12.8 jss = 2.17E-5
+ jsws = 8.200000000000001E-10 cjs = {7.433E-04*sw_func_psd_nw_cj} mjs = 0.34629
+ mjsws = 0.26859 cjsws = {9.2435E-11*sw_func_psd_nw_cj} cjswgs = {2.4701E-10*sw_func_psd_nw_cj}
+ mjswgs = 0.70393 pbs = 0.6587 pbsws = 0.7418
+ pbswgs = 1.3925 xrcrg1 = 12 xrcrg2 = 1
+ rbpb = 50 rbpd = 50 rbps = 50
+ rbdb = 50 rbsb = 50 gbmin = 1E-12
+ tnom = 30 ute = 5.591784564508111 lute = -6.91793810422675E-6
+ wute = -2.694665368921171E-6 pute = 2.822764647878656E-12 kt1 = 0.144080554246774
+ lkt1 = -6.884603388103184E-7 wkt1 = -3.028992661160058E-7 pkt1 = 3.369369883185032E-13
+ kt1l = 0 kt2 = -0.07901434332 lkt2 = 4.009909764692303E-8
+ wkt2 = 1.040075713246618E-8 pkt2 = -1.538838273731933E-14 ua1 = 7.80627001890499E-9
+ lua1 = -7.86960459150056E-15 wua1 = -2.512758996976034E-15 pua1 = 2.273923881335756E-21
+ ub1 = -1.209058997819079E-18 lub1 = 1.152961318315822E-24 wub1 = -2.116841066427713E-25
+ pub1 = 7.264328542281294E-31 uc1 = 2.661907042570155E-11 luc1 = -8.576043094614665E-17
+ wuc1 = -1.233837284487843E-17 puc1 = 8.010436116011549E-23 at = 1.77781670312476E5
+ lat = -0.091076202565067 wat = -0.079550045682395 pat = 6.128175602331857E-8
+ prt = 0 njs = 1.2556 xtis = 2
+ tpb = 1.9551E-3 tpbsw = 1.4242E-4 tpbswg = 0
+ tcj = 1.2407E-3 tcjsw = 0 tcjswg = 2E-12
+ tvoff = 0 tvfbsdoff = 0 saref = 3E-6
+ sbref = 3E-6 wlod = 0 ku0 = 4.5E-8
+ kvsat = 0.4 kvth0 = 2.65E-8 tku0 = 0
+ llodku0 = 0 wlodku0 = 1 llodvth = 0
+ wlodvth = 1 lku0 = 0 wku0 = 2.5E-7
+ pku0 = 0 lkvth0 = 0 wkvth0 = 2.5E-7
+ pkvth0 = 0 stk2 = 0 lodk2 = 1
+ steta0 = 0 lodeta0 = 1

.model phighvt_model.45 pmos
+ level = 54 lmin = 5E-7 lmax = 1E-6 wmin = 4.2E-7
+ wmax = 5.5E-7 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 4.23E-9
+ toxm = 4.23E-9 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 9.999999999999999E22 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {9.364E-9+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {-1.176E-8-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = -5.722E-9 dwb = -1.7864E-8 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = -1.002922590203037 lvth0 = -1.941857239753875E-9
+ wvth0 = -5.377182973878596E-8 pvth0 = 1.076235270137782E-14 k1 = 0.967674296935047
+ lk1 = -3.842320717088793E-7 wk1 = -2.035515704520215E-7 pk1 = 1.625267800725563E-13
+ k2 = -0.181390423301022 lk2 = 1.496523665746917E-7 wk2 = 7.76574175959613E-8
+ pk2 = -6.126170692025474E-14 k3 = -13.778 k3b = 2
+ w0 = 0 lpe0 = 0 lpeb = 0
+ vbm = -3 dvtp0 = 0 dvtp1 = 0
+ dvt0 = 4.05 dvt1 = 0.3 dvt2 = 0.03
+ dvt0w = -4.254 dvt1w = 1.1472E6 dvt2w = -8.96E-3
+ vfbsdoff = 0 u0 = -8.156766210691469E-3 lu0 = 1.311274477408242E-8
+ wu0 = 7.124172477522225E-9 pu0 = -6.039993490118817E-15 ua = -4.862971221307848E-9
+ lua = 3.40436989634035E-15 wua = 1.597918956113211E-15 pua = -1.513581819474104E-21
+ ub = 3.542203738837742E-18 lub = -2.184878095411868E-24 wub = -1.006902403662673E-24
+ pub = 9.67042959749419E-31 uc = 1.26565558777393E-10 luc = -1.413207068372154E-16
+ wuc = -8.775541556873272E-17 puc = 7.237678501124524E-23 ud = 0
+ up = 0 lp = 1 eu = 1.67
+ vsat = 1.412180674617322E5 lvsat = -0.054988313737967 wvsat = -0.072224272092402
+ pvsat = 5.45209030807453E-8 a0 = 1.334249587358845 la0 = 3.243962910533068E-7
+ wa0 = 3.858963040213183E-8 pa0 = -2.53720022141014E-13 ags = -1.663548076032844
+ lags = 1.525300688764714E-6 wags = 8.02131309738165E-7 pags = -4.199317832741241E-13
+ b0 = -3.801095781263752E-7 lb0 = 1.9899496634072E-13 wb0 = 9.99014260726699E-14
+ pb0 = -5.230039457756414E-20 b1 = -2.172690281833353E-9 lb1 = 1.137446816345397E-15
+ wb1 = 1.018652141859936E-15 pb1 = -5.332847693065135E-22 keta = 0.171044381795676
+ lketa = -1.355405130820674E-7 wketa = -6.778403675934686E-8 pketa = 4.781500184629057E-14
+ a1 = 0 a2 = 2.666671945779288 la2 = -1.910576069944018E-6
+ wa2 = -8.204683169563468E-7 pa2 = 8.3976573177116E-13 rdsw = 531.92
+ rdswmin = 0 rdw = 0 rdwmin = 0
+ rsw = 0 rswmin = 0 prwb = -0.32348
+ prwg = 0.02 wr = 1 voff = -0.282238518139819
+ lvoff = 3.883191231703363E-8 wvoff = 2.847266362559864E-8 pvoff = -1.365599153497132E-14
+ voffl = 0 minv = 0 nfactor = -4.460810936557472
+ lnfactor = 3.216959429887779E-6 wnfactor = 2.654039801880638E-6 pnfactor = -1.05765351637345E-12
+ eta0 = 4.257748279249928 leta0 = -3.003352813325579E-6 weta0 = -1.733675242928777E-6
+ peta0 = 1.321269412337004E-12 etab = 5.341684242148632 letab = -2.798607905663923E-6
+ wetab = -2.83868713540642E-6 petab = 1.486962633211878E-12 dsub = -7.58219479709538
+ ldsub = 5.688755996372296E-6 wdsub = 3.754703868431257E-6 pdsub = -2.600960483024024E-12
+ cit = 1E-5 cdsc = 0 cdscb = 0
+ cdscd = 0 pclm = 0.98956728602025 lpclm = 3.443778644645679E-7
+ wpclm = -8.32881057443681E-8 ppclm = -2.942915172258114E-13 pdiblc1 = 0.502671841132051
+ lpdiblc1 = -1.34733352692247E-7 wpdiblc1 = 1.120594246541181E-7 ppdiblc1 = -1.074604836970124E-13
+ pdiblc2 = -2.471606440192431E-3 lpdiblc2 = 2.969852223665756E-9 wpdiblc2 = 1.333705515404897E-9
+ ppdiblc2 = -1.36507426912722E-15 pdiblcb = 0.178684406608356 lpdiblcb = -4.131790638517839E-7
+ wpdiblcb = -2.144662220676342E-7 ppdiblcb = 2.19510467610665E-13 drout = 1.863642549847986
+ ldrout = -1.496250454558572E-6 wdrout = -4.740706527378017E-7 pdrout = 6.671601068084844E-13
+ pscbe1 = 3.631444187051065E9 lpscbe1 = -2.898039754330506E3 wpscbe1 = -1.136179271826355E3
+ ppscbe1 = 1.162902208299711E-3 pscbe2 = -2.856967350314064E-7 lpscbe2 = 3.020381081070891E-13
+ wpscbe2 = 1.182697201552993E-13 ppscbe2 = -1.211767958990995E-19 pvag = 0
+ delta = 0.01 fprout = 0 pdits = 0
+ pditsl = 0 pditsd = 0 lambda = 0
+ vtl = 0 lc = 5E-9 xn = 3
+ alpha0 = 2.45998434810948E-10 lalpha0 = -7.643310059222751E-17 walpha0 = -7.756488045888197E-17
+ palpha0 = 4.06067662178339E-23 alpha1 = 1.363722822892307E-9 lalpha1 = -6.615841722405806E-16
+ walpha1 = -6.713805515636419E-16 palpha1 = 3.514811463545978E-22 beta0 = 4.846188917724733
+ lbeta0 = 2.328559137759595E-6 wbeta0 = -2.32917110708429E-7 pbeta0 = -1.150195690359468E-13
+ aigbacc = 0.43 bigbacc = 0.054 cigbacc = 0.075
+ nigbacc = 1 aigbinv = 0.35 bigbinv = 0.03
+ cigbinv = 6E-3 eigbinv = 1.1 nigbinv = 3
+ aigc = 0.43 bigc = 0.054 cigc = 0.075
+ aigsd = 0.43 bigsd = 0.054 cigsd = 0.075
+ dlcig = 0 nigc = 1 poxedge = 1
+ pigcd = 1 ntox = 1 toxref = 4.23E-9
+ agidl = 2.735422469009476E-9 lagidl = -1.093201728972132E-15 wagidl = -6.192088945974723E-16
+ pagidl = 3.981929731310662E-22 bgidl = 1E9 cgidl = 300
+ egidl = 0.1 noia = 1.2E41 noib = 2E25
+ noic = 0 em = 4.1E7 af = 1
+ ef = 0.88 kf = 0 lintnoi = -6E-8
+ tnoia = 1.5 tnoib = 3.5 ntnoi = 1
+ rnoia = 0.577 rnoib = 0.37 xpart = 0
+ cgso = {5.932020000000001E-11/sw_func_tox_lv_ratio} cgdo = {5.932020000000001E-11/sw_func_tox_lv_ratio} cgbo = {0/sw_func_tox_lv_ratio}
+ ckappas = 0.6 cf = 1.2E-11 clc = 1E-7
+ cle = 0.6 dlc = -2.56E-9 dwc = 0
+ vfbcv = -0.1446893 noff = 4 voffcv = -0.1375
+ acde = 0.552 moin = 14.504 cgsl = {7.513892E-12/sw_func_tox_lv_ratio}
+ cgdl = {7.513892E-12/sw_func_tox_lv_ratio} ijthsrev = 0.1 ijthsfwd = 0.1
+ xjbvs = 1 bvs = 12.8 jss = 2.17E-5
+ jsws = 8.200000000000001E-10 cjs = {7.433E-04*sw_func_psd_nw_cj} mjs = 0.34629
+ mjsws = 0.26859 cjsws = {9.2435E-11*sw_func_psd_nw_cj} cjswgs = {2.4701E-10*sw_func_psd_nw_cj}
+ mjswgs = 0.70393 pbs = 0.6587 pbsws = 0.7418
+ pbswgs = 1.3925 xrcrg1 = 12 xrcrg2 = 1
+ rbpb = 50 rbpd = 50 rbps = 50
+ rbdb = 50 rbsb = 50 gbmin = 1E-12
+ tnom = 30 ute = -1.913212339972045 lute = 7.635763274467802E-7
+ wute = 9.250001751182367E-9 pute = 5.525318768808917E-14 kt1 = -0.639978433098398
+ lkt1 = 1.140397159172117E-7 wkt1 = 8.816749070110831E-8 pkt1 = -6.33276586189494E-14
+ kt1l = 0 kt2 = -0.019202376295926 lkt2 = -2.11196468415566E-8
+ wkt2 = -9.485999594195096E-9 pkt2 = 4.966110507553016E-15 ua1 = -2.614218264796126E-9
+ lua1 = 2.795973576633206E-15 wua1 = -5.730163198501746E-18 pua1 = -2.920702706122228E-22
+ ub1 = 9.592871998040652E-19 lub1 = -1.066384381875418E-24 wub1 = 9.020441011647798E-25
+ pub1 = -4.134902410270553E-31 uc1 = -4.651346300806516E-11 luc1 = -1.090782032601772E-17
+ wuc1 = 1.349515795718511E-16 puc1 = -7.064985093745546E-23 at = 9.80105852663166E4
+ lat = -9.428901598622055E-3 wat = -0.040278613467052 pat = 2.108665972227103E-8
+ prt = 0 njs = 1.2556 xtis = 2
+ tpb = 1.9551E-3 tpbsw = 1.4242E-4 tpbswg = 0
+ tcj = 1.2407E-3 tcjsw = 0 tcjswg = 2E-12
+ tvoff = 0 tvfbsdoff = 0 saref = 2.75E-6
+ sbref = 2.74E-6 wlod = 0 ku0 = 4.5E-8
+ kvsat = 0.4 kvth0 = 2.65E-8 tku0 = 0
+ llodku0 = 0 wlodku0 = 1 llodvth = 0
+ wlodvth = 1 lku0 = 0 wku0 = 2.5E-7
+ pku0 = 0 lkvth0 = 0 wkvth0 = 2.5E-7
+ pkvth0 = 0 stk2 = 0 lodk2 = 1
+ steta0 = 0 lodeta0 = 1

.model phighvt_model.46 pmos
+ level = 54 lmin = 2.5E-7 lmax = 5E-7 wmin = 4.2E-7
+ wmax = 5.5E-7 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 4.23E-9
+ toxm = 4.23E-9 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 9.999999999999999E22 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {9.364E-9+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {-1.176E-8-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = -5.722E-9 dwb = -1.7864E-8 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = -0.870589176251392 lvth0 = -7.122104611171923E-8
+ wvth0 = -1.054363305801525E-7 pvth0 = 3.780975218185004E-14 k1 = -0.442307409458575
+ lk1 = 3.539215512223094E-7 wk1 = 2.238538476380561E-7 pk1 = -6.122850440596109E-14
+ k2 = 0.298724166665139 lk2 = -1.016972235643927E-7 wk2 = -5.551445859767239E-8
+ pk2 = 8.45643370463636E-15 k3 = -13.778 k3b = 2
+ w0 = 0 lpe0 = 0 lpeb = 0
+ vbm = -3 dvtp0 = 0 dvtp1 = 0
+ dvt0 = 4.05 dvt1 = 0.3 dvt2 = 0.03
+ dvt0w = -4.254 dvt1w = 1.1472E6 dvt2w = -8.96E-3
+ vfbsdoff = 0 u0 = 0.033220659007765 lu0 = -8.549164876283849E-9
+ wu0 = -9.438744613659993E-9 pu0 = 2.631024865456899E-15 ua = 6.332939282885062E-9
+ lua = -2.456913170814722E-15 wua = -2.708157150278865E-15 pua = 7.407351437442752E-22
+ ub = -3.896037419134134E-18 lub = 1.709189915609568E-24 wub = 1.759637653535747E-24
+ pub = -4.812960909950972E-31 uc = -3.005267395215781E-10 luc = 8.227065316826204E-17
+ wuc = 1.057402794108092E-16 puc = -2.892208122444452E-23 ud = 0
+ up = 0 lp = 1 eu = 1.67
+ vsat = 2.43732056174395E5 lvsat = -0.10865643710882 wvsat = -0.073104381228718
+ pvsat = 5.498165781578907E-8 a0 = 2.815568624909638 la0 = -4.511038514852842E-7
+ wa0 = -9.340703153315596E-7 pa0 = 2.554869126494882E-13 ags = 1.25
+ b0 = 0 b1 = 0 keta = -0.15310787533246
+ lketa = 3.415967656965436E-8 wketa = 4.931481168814919E-8 pketa = -1.348858729294257E-14
+ a1 = 0 a2 = -2.553146660534578 la2 = 8.221033668334177E-7
+ wa2 = 1.640936633912694E-6 pa2 = -4.488289881077999E-13 rdsw = 531.92
+ rdswmin = 0 rdw = 0 rdwmin = 0
+ rsw = 0 rswmin = 0 prwb = -0.32348
+ prwg = 0.02 wr = 1 voff = -0.149909030180497
+ lvoff = -3.044522121943038E-8 wvoff = 5.000069305208339E-9 pvoff = -1.367618956360585E-15
+ voffl = 0 minv = 0 nfactor = 1.423107871092848
+ lnfactor = 1.366102557066842E-7 wnfactor = 1.327157602828407E-6 pnfactor = -3.630041475256258E-13
+ eta0 = -3.633444936690627 leta0 = 1.12784465908362E-6 weta0 = 1.654622996635722E-6
+ peta0 = -4.525724820398025E-13 etab = -8.510646857085425E-3 letab = 2.326122628350005E-9
+ wetab = 3.412576335636382E-9 petab = -9.33407879323263E-16 dsub = 6.15287208907249
+ ldsub = -1.501826219874307E-6 wdsub = -2.541191655291566E-6 pdsub = 6.95066741555349E-13
+ cit = 1E-5 cdsc = 0 cdscb = 0
+ cdscd = 0 pclm = 2.545313091341957 lpclm = -4.700861795374522E-7
+ wpclm = -1.351578025380412E-6 ppclm = 3.696836215020503E-13 pdiblc1 = 0.308268370164818
+ lpdiblc1 = -3.295924757148107E-8 wpdiblc1 = -1.951805348083544E-7 ppdiblc1 = 5.338577988078108E-14
+ pdiblc2 = -0.029055894063587 lpdiblc2 = 1.688725848026506E-8 wpdiblc2 = 8.742895882265783E-9
+ ppdiblc2 = -5.24393360998623E-15 pdiblcb = -1.032368813216711 lpdiblcb = 2.208315177910348E-7
+ wpdiblcb = 4.289324441352685E-7 ppdiblcb = -1.173216021198786E-13 drout = -3.174391179992618
+ ldrout = 1.141260963687581E-6 wdrout = 1.675898554748762E-6 pdrout = -4.583917726948813E-13
+ pscbe1 = -4.862853965286132E9 lpscbe1 = 1.548895214381062E3 wpscbe1 = 2.27235854365271E3
+ ppscbe1 = -6.215355088598892E-4 pscbe2 = 5.996865424990046E-7 lpscbe2 = -1.614777453456318E-13
+ wpscbe2 = -2.370409280135891E-13 ppscbe2 = 6.483543463027687E-20 pvag = 0
+ delta = 0.01 fprout = 0 pdits = 0
+ pditsl = 0 pditsd = 0 lambda = 0
+ vtl = 0 lc = 5E-9 xn = 3
+ alpha0 = 1E-10 alpha1 = 1E-10 beta0 = 9.52259235970739
+ lbeta0 = -1.19631592187166E-7 wbeta0 = -9.478253393360943E-7 pbeta0 = 2.592491868152085E-13
+ aigbacc = 0.43 bigbacc = 0.054 cigbacc = 0.075
+ nigbacc = 1 aigbinv = 0.35 bigbinv = 0.03
+ cigbinv = 6E-3 eigbinv = 1.1 nigbinv = 3
+ aigc = 0.43 bigc = 0.054 cigc = 0.075
+ aigsd = 0.43 bigsd = 0.054 cigsd = 0.075
+ dlcig = 0 nigc = 1 poxedge = 1
+ pigcd = 1 ntox = 1 toxref = 4.23E-9
+ agidl = 3.387373715009486E-9 lagidl = -1.434511245278057E-15 wagidl = -1.803984078321788E-15
+ pagidl = 1.01844647731442E-21 bgidl = 1E9 cgidl = 300
+ egidl = 0.1 noia = 1.2E41 noib = 2E25
+ noic = 0 em = 4.1E7 af = 1
+ ef = 0.88 kf = 0 lintnoi = -6E-8
+ tnoia = 1.5 tnoib = 3.5 ntnoi = 1
+ rnoia = 0.577 rnoib = 0.37 xpart = 0
+ cgso = {5.932020000000001E-11/sw_func_tox_lv_ratio} cgdo = {5.932020000000001E-11/sw_func_tox_lv_ratio} cgbo = {0/sw_func_tox_lv_ratio}
+ ckappas = 0.6 cf = 1.2E-11 clc = 1E-7
+ cle = 0.6 dlc = -2.56E-9 dwc = 0
+ vfbcv = -0.1446893 noff = 4 voffcv = -0.1375
+ acde = 0.552 moin = 14.504 cgsl = {7.513892E-12/sw_func_tox_lv_ratio}
+ cgdl = {7.513892E-12/sw_func_tox_lv_ratio} ijthsrev = 0.1 ijthsfwd = 0.1
+ xjbvs = 1 bvs = 12.8 jss = 2.17E-5
+ jsws = 8.200000000000001E-10 cjs = {7.433E-04*sw_func_psd_nw_cj} mjs = 0.34629
+ mjsws = 0.26859 cjsws = {9.2435E-11*sw_func_psd_nw_cj} cjswgs = {2.4701E-10*sw_func_psd_nw_cj}
+ mjswgs = 0.70393 pbs = 0.6587 pbsws = 0.7418
+ pbswgs = 1.3925 xrcrg1 = 12 xrcrg2 = 1
+ rbpb = 50 rbpd = 50 rbps = 50
+ rbdb = 50 rbsb = 50 gbmin = 1E-12
+ tnom = 30 ute = -2.577524172371553 lute = 1.111356857944571E-6
+ wute = 1.079212660132435E-6 pute = -5.048936632276642E-13 kt1 = -0.023707494793846
+ lkt1 = -2.085904457039871E-7 wkt1 = -1.763305400472213E-7 pkt1 = 7.514235043841608E-14
+ kt1l = 0 kt2 = -0.07837421088 lkt2 = 9.857991999897597E-9
+ ua1 = 5.388585636188553E-9 lua1 = -1.393654321610293E-15 wua1 = -1.18028050259961E-15
+ pua1 = 3.228303230710452E-22 ub1 = -2.316421710055975E-18 lub1 = 6.485147466145102E-25
+ wub1 = 2.349915472589213E-25 pub1 = -6.427488800626013E-32 uc1 = 2.059893257071996E-11
+ luc1 = -4.60425016594233E-17 wuc1 = -3.924840215773457E-17 puc1 = 2.05473234976172E-23
+ at = 1.8673869728E5 lat = -0.055879842800026 wat = -0.0538248422494
+ pat = 2.817838141440604E-8 prt = 0 njs = 1.2556
+ xtis = 2 tpb = 1.9551E-3 tpbsw = 1.4242E-4
+ tpbswg = 0 tcj = 1.2407E-3 tcjsw = 0
+ tcjswg = 2E-12 tvoff = 0 tvfbsdoff = 0
+ saref = 1.75E-6 sbref = 1.74E-6 wlod = 0
+ ku0 = 4.5E-8 kvsat = 0.4 kvth0 = 2.65E-8
+ tku0 = 0 llodku0 = 0 wlodku0 = 1
+ llodvth = 0 wlodvth = 1 lku0 = 0
+ wku0 = 2.5E-7 pku0 = 0 lkvth0 = 0
+ wkvth0 = 2.5E-7 pkvth0 = 0 stk2 = 0
+ lodk2 = 1 steta0 = 0 lodeta0 = 1

.model phighvt_model.47 pmos
+ level = 54 lmin = 1.8E-7 lmax = 2.5E-7 wmin = 4.2E-7
+ wmax = 5.5E-7 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 4.23E-9
+ toxm = 4.23E-9 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 9.999999999999999E22 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {9.364E-9+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {-1.176E-8-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = -5.722E-9 dwb = -1.7864E-8 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = -1.130976153846154 wvth0 = 3.279762738215387E-8
+ k1 = 0.85164386 k2 = -0.073084927969231 wk2 = -2.45974005959308E-8
+ k3 = -13.778 k3b = 2 w0 = 0
+ lpe0 = 0 lpeb = 0 vbm = -3
+ dvtp0 = 0 dvtp1 = 0 dvt0 = 4.05
+ dvt1 = 0.3 dvt2 = 0.03 dvt0w = -4.254
+ dvt1w = 1.1472E6 dvt2w = -8.96E-3 vfbsdoff = 0
+ u0 = 2.836800725274724E-3 lu0 = -2.38571958857143E-10 wu0 = 1.803869506018466E-10
+ ua = -2.649633E-9 ub = 2.3528289E-18 uc = 2.58041E-13
+ ud = 0 up = 0 lp = 1
+ eu = 1.67 vsat = -1.535201999999999E5 wvsat = 0.1279107467904
+ a0 = 1.166315 ags = 1.25 b0 = 0
+ b1 = 0 keta = -0.028218739 a1 = 0
+ a2 = 0.45249595 rdsw = 531.92 rdswmin = 0
+ rdw = 0 rdwmin = 0 rsw = 0
+ rswmin = 0 prwb = -0.32348 prwg = 0.02
+ wr = 1 voff = -0.26121797 voffl = 0
+ minv = 0 nfactor = 1.9225604 eta0 = 0.49
+ etab = -6.25E-6 dsub = 0.66213569 cit = 1E-5
+ cdsc = 0 cdscb = 0 cdscd = 0
+ pclm = 0.82665932 pdiblc1 = 0.18776805 pdiblc2 = 0.03268459467678
+ wpdiblc2 = -1.042913398752886E-8 pdiblcb = -0.225 drout = 0.9981043
+ pscbe1 = 7.9996855E8 pscbe2 = 9.3174823E-9 pvag = 0
+ delta = 0.01 fprout = 0 pdits = 0
+ pditsl = 0 pditsd = 0 lambda = 0
+ vtl = 0 lc = 5E-9 xn = 3
+ alpha0 = 1E-10 alpha1 = 1E-10 beta0 = 9.0852145
+ aigbacc = 0.43 bigbacc = 0.054 cigbacc = 0.075
+ nigbacc = 1 aigbinv = 0.35 bigbinv = 0.03
+ cigbinv = 6E-3 eigbinv = 1.1 nigbinv = 3
+ aigc = 0.43 bigc = 0.054 cigc = 0.075
+ aigsd = 0.43 bigsd = 0.054 cigsd = 0.075
+ dlcig = 0 nigc = 1 poxedge = 1
+ pigcd = 1 ntox = 1 toxref = 4.23E-9
+ agidl = -1.857256459303387E-9 wagidl = 1.919496754211189E-15 bgidl = 1E9
+ cgidl = 300 egidl = 0.1 noia = 1.2E41
+ noib = 2E25 noic = 0 em = 4.1E7
+ af = 1 ef = 0.88 kf = 0
+ lintnoi = -6E-8 tnoia = 1.5 tnoib = 3.5
+ ntnoi = 1 rnoia = 0.577 rnoib = 0.37
+ xpart = 0 cgso = {5.932020000000001E-11/sw_func_tox_lv_ratio} cgdo = {5.932020000000001E-11/sw_func_tox_lv_ratio}
+ cgbo = {0/sw_func_tox_lv_ratio} ckappas = 0.6 cf = 1.2E-11
+ clc = 1E-7 cle = 0.6 dlc = -2.56E-9
+ dwc = 0 vfbcv = -0.1446893 noff = 4
+ voffcv = -0.1375 acde = 0.552 moin = 14.504
+ cgsl = {7.513892E-12/sw_func_tox_lv_ratio} cgdl = {7.513892E-12/sw_func_tox_lv_ratio} ijthsrev = 0.1
+ ijthsfwd = 0.1 xjbvs = 1 bvs = 12.8
+ jss = 2.17E-5 jsws = 8.200000000000001E-10 cjs = {7.433E-04*sw_func_psd_nw_cj}
+ mjs = 0.34629 mjsws = 0.26859 cjsws = {9.2435E-11*sw_func_psd_nw_cj}
+ cjswgs = {2.4701E-10*sw_func_psd_nw_cj} mjswgs = 0.70393 pbs = 0.6587
+ pbsws = 0.7418 pbswgs = 1.3925 xrcrg1 = 12
+ xrcrg2 = 1 rbpb = 50 rbpd = 50
+ rbps = 50 rbdb = 50 rbsb = 50
+ gbmin = 1E-12 tnom = 30 ute = 1.485640707507692
+ wute = -7.666986561430265E-7 kt1 = -0.786322461538461 wkt1 = 9.839288214646141E-8
+ kt1l = 0 kt2 = -0.042333 ua1 = 2.9333E-10
+ ub1 = 5.4574E-20 uc1 = -1.477342849615384E-10 wuc1 = 3.587342987508644E-17
+ at = -1.756023076923074E4 wat = 0.049196441073231 prt = 0
+ njs = 1.2556 xtis = 2 tpb = 1.9551E-3
+ tpbsw = 1.4242E-4 tpbswg = 0 tcj = 1.2407E-3
+ tcjsw = 0 tcjswg = 2E-12 tvoff = 0
+ tvfbsdoff = 0 saref = 1.1E-6 sbref = 1.1E-6
+ wlod = 0 ku0 = 4.5E-8 kvsat = 0.4
+ kvth0 = 2.65E-8 tku0 = 0 llodku0 = 0
+ wlodku0 = 1 llodvth = 0 wlodvth = 1
+ lku0 = 0 wku0 = 2.5E-7 pku0 = 0
+ lkvth0 = 0 wkvth0 = 2.5E-7 pkvth0 = 0
+ stk2 = 0 lodk2 = 1 steta0 = 0
+ lodeta0 = 1

.model phighvt_model.48 pmos
+ level = 54 lmin = 1.5E-7 lmax = 1.8E-7 wmin = 4.2E-7
+ wmax = 5.5E-7 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 4.23E-9
+ toxm = 4.23E-9 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 9.999999999999999E22 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {9.364E-9+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {-1.176E-8-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = -5.722E-9 dwb = -1.7864E-8 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = -1.488046499692308 lvth0 = 7.267095678660915E-8
+ wvth0 = 2.224991041605315E-7 pvth0 = -3.860804455393541E-14 k1 = 0.85164386
+ k2 = -0.073084927969231 wk2 = -2.45974005959308E-8 k3 = -13.778
+ k3b = 2 w0 = 0 lpe0 = 0
+ lpeb = 0 vbm = -3 dvtp0 = 0
+ dvtp1 = 0 dvt0 = 4.05 dvt1 = 0.3
+ dvt2 = 0.03 dvt0w = -4.254 dvt1w = 1.1472E6
+ dvt2w = -8.96E-3 vfbsdoff = 0 u0 = 2.28576663507692E-3
+ lu0 = -1.264255008200858E-10 wu0 = 4.649391657694135E-10 pu0 = -5.791206683090322E-17
+ ua = -2.649633E-9 ub = 2.3528289E-18 uc = 2.58041E-13
+ ud = 0 up = 0 lp = 1
+ eu = 1.67 vsat = -1.367559375876921E6 lvsat = 0.247081253074471
+ wvsat = 0.772895767836883 pvsat = -1.312673514833803E-7 a0 = 1.166315
+ ags = 1.25 b0 = 0 b1 = 0
+ keta = -0.028218739 a1 = 0 a2 = 0.45249595
+ rdsw = 531.92 rdswmin = 0 rdw = 0
+ rdwmin = 0 rsw = 0 rswmin = 0
+ prwb = -0.32348 prwg = 0.02 wr = 1
+ voff = -0.26121797 voffl = 0 minv = 0
+ nfactor = 1.9225604 eta0 = 0.49 etab = -6.25E-6
+ dsub = 0.66213569 cit = 1E-5 cdsc = 0
+ cdscb = 0 cdscd = 0 pclm = 0.82665932
+ pdiblc1 = 0.18776805 pdiblc2 = 0.03268459467678 wpdiblc2 = -1.042913398752886E-8
+ pdiblcb = -0.225 drout = 0.9981043 pscbe1 = 7.9996855E8
+ pscbe2 = 9.3174823E-9 pvag = 0 delta = 0.01
+ fprout = 0 pdits = 0 pditsl = 0
+ pditsd = 0 lambda = 0 vtl = 0
+ lc = 5E-9 xn = 3 alpha0 = 1E-10
+ alpha1 = 1E-10 beta0 = 9.0852145 aigbacc = 0.43
+ bigbacc = 0.054 cigbacc = 0.075 nigbacc = 1
+ aigbinv = 0.35 bigbinv = 0.03 cigbinv = 6E-3
+ eigbinv = 1.1 nigbinv = 3 aigc = 0.43
+ bigc = 0.054 cigc = 0.075 aigsd = 0.43
+ bigsd = 0.054 cigsd = 0.075 dlcig = 0
+ nigc = 1 poxedge = 1 pigcd = 1
+ ntox = 1 toxref = 4.23E-9 agidl = 1.120381351327833E-8
+ lagidl = -2.658188960819832E-15 wagidl = -5.019484012262248E-15 pagidl = 1.412221365592674E-21
+ bgidl = 1E9 cgidl = 300 egidl = 0.1
+ noia = 1.2E41 noib = 2E25 noic = 0
+ em = 4.1E7 af = 1 ef = 0.88
+ kf = 0 lintnoi = -6E-8 tnoia = 1.5
+ tnoib = 3.5 ntnoi = 1 rnoia = 0.577
+ rnoib = 0.37 xpart = 0 cgso = {5.932020000000001E-11/sw_func_tox_lv_ratio}
+ cgdo = {5.932020000000001E-11/sw_func_tox_lv_ratio} cgbo = {0/sw_func_tox_lv_ratio} ckappas = 0.6
+ cf = 1.2E-11 clc = 1E-7 cle = 0.6
+ dlc = -2.56E-9 dwc = 0 vfbcv = -0.1446893
+ noff = 4 voffcv = -0.1375 acde = 0.552
+ moin = 14.504 cgsl = {7.513892E-12/sw_func_tox_lv_ratio} cgdl = {7.513892E-12/sw_func_tox_lv_ratio}
+ ijthsrev = 0.1 ijthsfwd = 0.1 xjbvs = 1
+ bvs = 12.8 jss = 2.17E-5 jsws = 8.200000000000001E-10
+ cjs = {7.433E-04*sw_func_psd_nw_cj} mjs = 0.34629 mjsws = 0.26859
+ cjsws = {9.2435E-11*sw_func_psd_nw_cj} cjswgs = {2.4701E-10*sw_func_psd_nw_cj} mjswgs = 0.70393
+ pbs = 0.6587 pbsws = 0.7418 pbswgs = 1.3925
+ xrcrg1 = 12 xrcrg2 = 1 rbpb = 50
+ rbpd = 50 rbps = 50 rbdb = 50
+ rbsb = 50 gbmin = 1E-12 tnom = 30
+ ute = 10.792456103021516 lute = -1.894123069294974E-6 wute = -5.711149084948447E-6
+ pute = 1.00629455127048E-12 kt1 = -0.786322461538461 wkt1 = 9.839288214646141E-8
+ kt1l = 0 kt2 = -0.042333 ua1 = 2.9333E-10
+ ub1 = 1.839925729230766E-18 lub1 = -3.633547839330455E-25 wub1 = -9.485073838918873E-25
+ pub1 = 1.930402227696769E-31 uc1 = -1.477342849615384E-10 wuc1 = 3.587342987508644E-17
+ at = -9.102360953846134E5 lat = 0.181677391966523 wat = 0.523450133019174
+ pat = -9.652011138483845E-8 prt = 0 njs = 1.2556
+ xtis = 2 tpb = 1.9551E-3 tpbsw = 1.4242E-4
+ tpbswg = 0 tcj = 1.2407E-3 tcjsw = 0
+ tcjswg = 2E-12 tvoff = 0 tvfbsdoff = 0
+ saref = 1.1E-6 sbref = 1.1E-6 wlod = 0
+ ku0 = 4.5E-8 kvsat = 0.4 kvth0 = 2.65E-8
+ tku0 = 0 llodku0 = 0 wlodku0 = 1
+ llodvth = 0 wlodvth = 1 lku0 = 0
+ wku0 = 2.5E-7 pku0 = 0 lkvth0 = 0
+ wkvth0 = 2.5E-7 pkvth0 = 0 stk2 = 0
+ lodk2 = 1 steta0 = 0 lodeta0 = 1

.ends sky130_fd_pr__pfet_01v8_hvt
