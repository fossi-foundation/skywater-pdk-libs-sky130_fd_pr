* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

******************************************************************
******************************************************************
*  *****************************************************
*  04/14/2021 Usman Suriono
*      Why     : New scalable sky130_fd_pr__nfet_01v8 native 5v model
*      What    : Converted from discrete nhvnative model
*      What    : Converted from discrete nshort model
*                Replaced rsh from 1 to calculated rsh from the original model.
*                PDK netlist nrd/nrs = ratio of distance the middle of the contact to Gate.
*
*  *****************************************************
*
*  Nmos Native 5V Model
*  -----------------------------------------------------

.subckt  sky130_fd_pr__nfet_05v0_nvt  d g s b  mult=1
+ 
.param  l = 1 w = 1 nf = 1 ad = 0 as = 0 pd = 0 ps = 0 nrd = {0.14/w} nrs = {0.14/w}
+ sa = 0 sb = 0 sd = 0
+ swx_nrds = {89.1*nf/w+443.5}

Msky130_fd_pr__nfet_05v0_nvt  d g s b nhvnative_model l = {l} w = {w} ad = {ad} as = {as} pd = {pd} ps = {ps} nrd = {nrd} nrs = {nrs} sa = {sa} sb = {sb} sd = {sd} nf = {nf}
* + deltox = 0.3*(sw_tox_hv_corner - sw_tox_hv_nom) + sw_tox_hv_mc + sw_mm_tox_hv * mismatch_factor*MC_MM_SWITCH*AGAUSS(0,1.0,1)/sqrt(l*w*mult)
* + mulu0  = sw_u0_sky130_fd_pr__nfet_01v8_nat**(0.17*10/w+0.83)
+ delvto = {sw_vth0_sky130_fd_pr__nfet_01v8_nat*(0.07*4/l+0.930)*(0.010*10/w+0.990)*(0.001*40/(w*l)+0.999)+sw_mm_vth0_sky130_fd_pr__nfet_01v8_nat*mismatch_factor*MC_MM_SWITCH*AGAUSS(0,1.0,1)/sqrt(l*w*mult)+sw_vth0_sky130_fd_pr__nfet_01v8_nat_mc*2}



.model nhvnative_model.1 nmos
+ level = 54 lmin = 8E-6 lmax = 2.525E-5 wmin = 1E-5
+ wmax = 1.01E-4 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 1.16E-8
+ toxm = 1.16E-8 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 1E23 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {4.5E-8+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {6.93E-8-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = -4.6E-9 dwb = 1.92E-9 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = 0.038459 lvth0 = 2.72244E-8
+ k1 = 0.364 k2 = 0.041446 lk2 = -1.271545E-8
+ k3 = 1.4 k3b = -0.58 w0 = 0
+ lpe0 = -1.236227E-14 lpeb = 0 vbm = -3
+ dvtp0 = 0 dvtp1 = 0 dvt0 = 5.7
+ dvt1 = 0.21851 dvt2 = 0.04 dvt0w = 7.7
+ dvt1w = 1.272E6 dvt2w = -0.032 vfbsdoff = 0
+ u0 = 4.45181E-2 lu0 = -2.145301E-9 ua = 1.096856E-9
+ lua = -2.413176E-17 ub = -1.500717E-19 lub = -1.033446E-24
+ uc = 1.9159E-11 ud = 0 up = 0
+ lp = 1 eu = 1.67 vsat = 7.5917E4
+ a0 = 1.387857 la0 = -1.035676E-5 ags = 2.90552E-2
+ lags = 3.780528E-6 b0 = 5.734E-8 b1 = 4.9905E-8
+ keta = -7.522213E-3 lketa = -1.067247E-7 a1 = 0
+ a2 = 0.962934 rdsw = 430 rdswmin = 0
+ rdw = 0 rdwmin = 0 rsw = 0
+ rswmin = 0 prwb = 0 prwg = 1E-12
+ wr = 1 voff = 0 voffl = 1.944533E-8
+ minv = 0 nfactor = 0.701166 lnfactor = -9.975764E-8
+ eta0 = 9 etab = -2.1692E-4 dsub = 0.42
+ cit = 9.258412E-8 cdsc = 0 cdscb = 1.415095E-7
+ cdscd = 1.5E-5 pclm = 0.089 pdiblc1 = 1.0772E-6
+ pdiblc2 = 5.1E-4 pdiblcb = 0 drout = 0.11135
+ pscbe1 = 2.7814E8 pscbe2 = 1.6E-8 pvag = 4.541944
+ delta = 7E-3 fprout = 0 pdits = -2.630332E-3
+ lpdits = 6.539373E-8 pditsl = 0 pditsd = 0
+ lambda = 0 vtl = 0 lc = 5E-9
+ xn = 3 alpha0 = 2.97923E-6 lalpha0 = -2.08346E-11
+ alpha1 = 0.5456 beta0 = 20.117451 lbeta0 = -8.73756E-6
+ aigbacc = 1 bigbacc = 0 cigbacc = 0
+ nigbacc = 1 aigbinv = 0.35 bigbinv = 0.03
+ cigbinv = 6E-3 eigbinv = 1.1 nigbinv = 3
+ aigc = 0.43 bigc = 0.054 cigc = 0.075
+ aigsd = 0.43 bigsd = 0.054 cigsd = 0.075
+ dlcig = 0 nigc = 1 poxedge = 1
+ pigcd = 1 ntox = 1 toxref = 1.16E-8
+ agidl = 0 bgidl = 2.3E9 cgidl = 0.5
+ egidl = 0.8 noia = 2.5E41 noib = 0
+ noic = 0 em = 4.1E7 af = 1
+ ef = 1 kf = 0 lintnoi = 0
+ tnoia = 7.6E6 tnoib = 7.2E6 ntnoi = 1
+ rnoia = 0.8 rnoib = 0.38 xpart = 0
+ cgso = {2.678273E-10/sw_func_tox_hv_ratio} cgdo = {2.678273E-10/sw_func_tox_hv_ratio} cgbo = {0/sw_func_tox_hv_ratio}
+ ckappas = 0.6 cf = 0 clc = 1E-7
+ cle = 0.6 dlc = 6.0712E-8 dwc = 0
+ vfbcv = -1 noff = 4 voffcv = 0.216
+ acde = 1.16 moin = 15 cgsl = {3.85585E-11/sw_func_tox_hv_ratio}
+ cgdl = {3.85585E-11/sw_func_tox_hv_ratio} ijthsrev = 0.1 ijthsfwd = 0.1
+ xjbvs = 1 bvs = 12.69 jss = 4.2966E-4
+ jsws = 8.04E-10 cjs = {8.310E-04*sw_func_nsd_pw_cj} mjs = 0.28329
+ mjsws = 0.057926 cjsws = {8.887314E-11*sw_func_nsd_pw_cj} cjswgs = {3.736446E-11*sw_func_nsd_pw_cj}
+ mjswgs = 0.33 pbs = 0.66345 pbsws = 1
+ pbswgs = 0.2442 xrcrg1 = 12 xrcrg2 = 1
+ rbpb = 50 rbpd = 50 rbps = 50
+ rbdb = 50 rbsb = 50 gbmin = 1E-12
+ tnom = 30 ute = -1.464 kt1 = -0.370524
+ lkt1 = 1.149679E-7 kt1l = 0 kt2 = -0.01144
+ ua1 = 1E-9 ub1 = -1.088076E-18 lub1 = 2.950191E-24
+ uc1 = 1E-11 at = 8.63772E4 lat = -0.496661
+ prt = 0 njs = 1.5764 xtis = 0
+ tpb = 1.9685E-3 tpbsw = 1E-3 tpbswg = 0
+ tcj = 8.3E-4 tcjsw = 0 tcjswg = 0
+ tvoff = 0 tvfbsdoff = 0 saref = 3E-6
+ sbref = 3E-6 wlod = 0 ku0 = -3E-8
+ kvsat = 0.4 kvth0 = -7E-9 tku0 = 0
+ llodku0 = 0 wlodku0 = 1 llodvth = 0
+ wlodvth = 1 lku0 = 0 wku0 = 2E-7
+ pku0 = 0 lkvth0 = 0 wkvth0 = 8E-7
+ pkvth0 = 0 stk2 = 0 lodk2 = 1
+ steta0 = 0 lodeta0 = 1

.model nhvnative_model.2 nmos
+ level = 54 lmin = 4E-6 lmax = 8E-6 wmin = 1E-5
+ wmax = 1.01E-4 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 1.16E-8
+ toxm = 1.16E-8 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 1E23 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {4.5E-8+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {6.93E-8-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = -4.6E-9 dwb = 1.92E-9 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = 2.65944E-2 lvth0 = 1.204967E-7
+ k1 = 0.364 k2 = 4.01426E-2 lk2 = -2.469461E-9
+ k3 = 1.4 k3b = -0.58 w0 = 0
+ lpe0 = -1.236227E-14 lpeb = 0 vbm = -3
+ dvtp0 = 0 dvtp1 = 0 dvt0 = 5.7
+ dvt1 = 0.21851 dvt2 = 0.04 dvt0w = 7.7
+ dvt1w = 1.272E6 dvt2w = -0.032 vfbsdoff = 0
+ u0 = 4.57121E-2 lu0 = -1.153225E-8 ua = 1.361378E-9
+ lua = -2.103649E-15 ub = -5.413346E-19 lub = 2.042428E-24
+ uc = 8.716809E-12 luc = 8.209024E-17 ud = 0
+ up = 0 lp = 1 eu = 1.67
+ vsat = 7.865956E4 lvsat = -2.15604E-2 a0 = 5.85431E-2
+ la0 = 9.350289E-8 ags = 0.323215 lags = 1.468017E-6
+ b0 = -2.154583E-7 lb0 = 2.144576E-12 b1 = 9.808079E-8
+ lb1 = -3.787292E-13 keta = -2.22506E-2 lketa = 9.061269E-9
+ a1 = 0 a2 = 0.962934 rdsw = 430
+ rdswmin = 0 rdw = 0 rdwmin = 0
+ rsw = 0 rswmin = 0 prwb = 0
+ prwg = 1E-12 wr = 1 voff = 0
+ voffl = 1.944533E-8 minv = 0 nfactor = 0.71299
+ lnfactor = -1.927151E-7 eta0 = 9 etab = -2.1692E-4
+ dsub = 0.42 cit = 9.258412E-8 cdsc = 0
+ cdscb = 1.415095E-7 cdscd = 1.5E-5 pclm = 6.15068E-2
+ lpclm = 2.161348E-7 pdiblc1 = 1.264381E-6 lpdiblc1 = -1.471508E-12
+ pdiblc2 = 8.092585E-4 lpdiblc2 = -2.352591E-9 pdiblcb = 0
+ drout = 9.20044E-2 ldrout = 1.520836E-7 pscbe1 = 3.103634E8
+ lpscbe1 = -253.320903 pscbe2 = 2.773866E-8 lpscbe2 = -9.228227E-14
+ pvag = 4.541944 delta = 7E-3 fprout = 0
+ pdits = 4.614531E-3 lpdits = 8.438971E-9 pditsl = 0
+ pditsd = 0 lambda = 0 vtl = 0
+ lc = 5E-9 xn = 3 alpha0 = -1.293773E-6
+ lalpha0 = 1.275719E-11 alpha1 = 0.981907 lalpha1 = -3.429986E-6
+ beta0 = 18.579315 lbeta0 = 3.354339E-6 aigbacc = 1
+ bigbacc = 0 cigbacc = 0 nigbacc = 1
+ aigbinv = 0.35 bigbinv = 0.03 cigbinv = 6E-3
+ eigbinv = 1.1 nigbinv = 3 aigc = 0.43
+ bigc = 0.054 cigc = 0.075 aigsd = 0.43
+ bigsd = 0.054 cigsd = 0.075 dlcig = 0
+ nigc = 1 poxedge = 1 pigcd = 1
+ ntox = 1 toxref = 1.16E-8 agidl = 0
+ bgidl = 2.3E9 cgidl = 0.5 egidl = 0.8
+ noia = 2.5E41 noib = 0 noic = 0
+ em = 4.1E7 af = 1 ef = 1
+ kf = 0 lintnoi = 0 tnoia = 7.6E6
+ tnoib = 7.2E6 ntnoi = 1 rnoia = 0.8
+ rnoib = 0.38 xpart = 0 cgso = {2.678273E-10/sw_func_tox_hv_ratio}
+ cgdo = {2.678273E-10/sw_func_tox_hv_ratio} cgbo = {0/sw_func_tox_hv_ratio} ckappas = 0.6
+ cf = 0 clc = 1E-7 cle = 0.6
+ dlc = 6.0712E-8 dwc = 0 vfbcv = -1
+ noff = 4 voffcv = 0.216 acde = 1.16
+ moin = 15 cgsl = {3.85585E-11/sw_func_tox_hv_ratio} cgdl = {3.85585E-11/sw_func_tox_hv_ratio}
+ ijthsrev = 0.1 ijthsfwd = 0.1 xjbvs = 1
+ bvs = 12.69 jss = 4.2966E-4 jsws = 8.04E-10
+ cjs = {8.310E-04*sw_func_nsd_pw_cj} mjs = 0.28329 mjsws = 0.057926
+ cjsws = {8.887314E-11*sw_func_nsd_pw_cj} cjswgs = {3.736446E-11*sw_func_nsd_pw_cj} mjswgs = 0.33
+ pbs = 0.66345 pbsws = 1 pbswgs = 0.2442
+ xrcrg1 = 12 xrcrg2 = 1 rbpb = 50
+ rbpd = 50 rbps = 50 rbdb = 50
+ rbsb = 50 gbmin = 1E-12 tnom = 30
+ ute = -1.153061 lute = -2.444418E-6 kt1 = -0.353313
+ lkt1 = -2.033853E-8 kt1l = 0 kt2 = -7.022558E-3
+ lkt2 = -3.472728E-8 ua1 = 1.540596E-9 lua1 = -4.249841E-15
+ ub1 = 1.679853E-19 lub1 = -6.924206E-24 uc1 = 5.768829E-11
+ luc1 = -3.748967E-16 at = 2.358614E4 lat = -3.035601E-3
+ prt = 0 njs = 1.5764 xtis = 0
+ tpb = 1.9685E-3 tpbsw = 1E-3 tpbswg = 0
+ tcj = 8.3E-4 tcjsw = 0 tcjswg = 0
+ tvoff = 0 tvfbsdoff = 0 saref = 3E-6
+ sbref = 3E-6 wlod = 0 ku0 = -3E-8
+ kvsat = 0.4 kvth0 = -7E-9 tku0 = 0
+ llodku0 = 0 wlodku0 = 1 llodvth = 0
+ wlodvth = 1 lku0 = 0 wku0 = 2E-7
+ pku0 = 0 lkvth0 = 0 wkvth0 = 8E-7
+ pkvth0 = 0 stk2 = 0 lodk2 = 1
+ steta0 = 0 lodeta0 = 1

.model nhvnative_model.3 nmos
+ level = 54 lmin = 2E-6 lmax = 4E-6 wmin = 1E-5
+ wmax = 1.01E-4 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 1.16E-8
+ toxm = 1.16E-8 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 1E23 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {4.5E-8+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {6.93E-8-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = -4.6E-9 dwb = 1.92E-9 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = 6.65513E-2 lvth0 = -3.379291E-8
+ k1 = 0.364 k2 = 4.03809E-2 lk2 = -3.389605E-9
+ k3 = 1.4 k3b = -0.58 w0 = 0
+ lpe0 = -1.236227E-14 lpeb = 0 vbm = -3
+ dvtp0 = 0 dvtp1 = 0 dvt0 = 5.7
+ dvt1 = 0.21851 dvt2 = 0.04 dvt0w = 7.7
+ dvt1w = 1.272E6 dvt2w = -0.032 vfbsdoff = 0
+ u0 = 4.25045E-2 lu0 = 8.538881E-10 ua = 8.189707E-10
+ lua = -9.196547E-18 ub = 5.293514E-20 lub = -2.522851E-25
+ uc = 2.754967E-11 luc = 9.36905E-18 ud = 0
+ up = 0 lp = 1 eu = 1.67
+ vsat = 7.692538E4 lvsat = -0.014864 a0 = 7.93386E-2
+ la0 = 1.320303E-8 ags = 0.538755 lags = 6.357341E-7
+ b0 = 3.3993E-7 b1 = 0 keta = -0.019904
+ a1 = 0 a2 = 0.962934 rdsw = 430
+ rdswmin = 0 rdw = 0 rdwmin = 0
+ rsw = 0 rswmin = 0 prwb = 0
+ prwg = 1E-12 wr = 1 voff = 0
+ voffl = 1.944533E-8 minv = 0 nfactor = 0.681365
+ lnfactor = -7.059671E-8 eta0 = 9 etab = -2.1692E-4
+ dsub = 0.42 cit = 9.258412E-8 cdsc = 0
+ cdscb = 1.415095E-7 cdscd = 1.5E-5 pclm = 0.11748
+ pdiblc1 = 8.833E-7 pdiblc2 = 2E-4 pdiblcb = 0
+ drout = 0.13139 pscbe1 = 2.4476E8 pscbe2 = 3.84E-9
+ pvag = 4.541944 delta = 7E-3 fprout = 0
+ pdits = -5.48524E-3 lpdits = 4.743823E-8 pditsl = 0
+ pditsd = 0 lambda = 0 vtl = 0
+ lc = 5E-9 xn = 3 alpha0 = 1.997342E-6
+ lalpha0 = 4.887575E-14 alpha1 = 0.093632 beta0 = 16.979784
+ lbeta0 = 9.530771E-6 aigbacc = 1 bigbacc = 0
+ cigbacc = 0 nigbacc = 1 aigbinv = 0.35
+ bigbinv = 0.03 cigbinv = 6E-3 eigbinv = 1.1
+ nigbinv = 3 aigc = 0.43 bigc = 0.054
+ cigc = 0.075 aigsd = 0.43 bigsd = 0.054
+ cigsd = 0.075 dlcig = 0 nigc = 1
+ poxedge = 1 pigcd = 1 ntox = 1
+ toxref = 1.16E-8 agidl = 0 bgidl = 2.3E9
+ cgidl = 0.5 egidl = 0.8 noia = 2.5E41
+ noib = 0 noic = 0 em = 4.1E7
+ af = 1 ef = 1 kf = 0
+ lintnoi = 0 tnoia = 7.6E6 tnoib = 7.2E6
+ ntnoi = 1 rnoia = 0.8 rnoib = 0.38
+ xpart = 0 cgso = {2.678273E-10/sw_func_tox_hv_ratio} cgdo = {2.678273E-10/sw_func_tox_hv_ratio}
+ cgbo = {0/sw_func_tox_hv_ratio} ckappas = 0.6 cf = 0
+ clc = 1E-7 cle = 0.6 dlc = 6.0712E-8
+ dwc = 0 vfbcv = -1 noff = 4
+ voffcv = 0.216 acde = 1.16 moin = 15
+ cgsl = {3.85585E-11/sw_func_tox_hv_ratio} cgdl = {3.85585E-11/sw_func_tox_hv_ratio} ijthsrev = 0.1
+ ijthsfwd = 0.1 xjbvs = 1 bvs = 12.69
+ jss = 4.2966E-4 jsws = 8.04E-10 cjs = {8.310E-04*sw_func_nsd_pw_cj}
+ mjs = 0.28329 mjsws = 0.057926 cjsws = {8.887314E-11*sw_func_nsd_pw_cj}
+ cjswgs = {3.736446E-11*sw_func_nsd_pw_cj} mjswgs = 0.33 pbs = 0.66345
+ pbsws = 1 pbswgs = 0.2442 xrcrg1 = 12
+ xrcrg2 = 1 rbpb = 50 rbpd = 50
+ rbps = 50 rbdb = 50 rbsb = 50
+ gbmin = 1E-12 tnom = 30 ute = -1.7861
+ kt1 = -0.35858 kt1l = 0 kt2 = -0.016016
+ ua1 = 4.4E-10 ub1 = -1.810968E-18 lub1 = 7.173235E-25
+ uc1 = -3.94E-11 at = 3.322384E4 lat = -4.02506E-2
+ prt = 0 njs = 1.5764 xtis = 0
+ tpb = 1.9685E-3 tpbsw = 1E-3 tpbswg = 0
+ tcj = 8.3E-4 tcjsw = 0 tcjswg = 0
+ tvoff = 0 tvfbsdoff = 0 saref = 3E-6
+ sbref = 3E-6 wlod = 0 ku0 = -3E-8
+ kvsat = 0.4 kvth0 = -7E-9 tku0 = 0
+ llodku0 = 0 wlodku0 = 1 llodvth = 0
+ wlodvth = 1 lku0 = 0 wku0 = 2E-7
+ pku0 = 0 lkvth0 = 0 wkvth0 = 8E-7
+ pkvth0 = 0 stk2 = 0 lodk2 = 1
+ steta0 = 0 lodeta0 = 1

.model nhvnative_model.4 nmos
+ level = 54 lmin = 1E-6 lmax = 2E-6 wmin = 1E-5
+ wmax = 1.01E-4 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 1.16E-8
+ toxm = 1.16E-8 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 1E23 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {4.5E-8+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {6.93E-8-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = -4.6E-9 dwb = 1.92E-9 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = 3.77066E-2 lvth0 = 1.989864E-8
+ k1 = 0.364 k2 = 3.69676E-2 lk2 = 2.964032E-9
+ k3 = 1.4 k3b = -0.58 w0 = 0
+ lpe0 = -1.236227E-14 lpeb = 0 vbm = -3
+ dvtp0 = 0 dvtp1 = 0 dvt0 = 5.7
+ dvt1 = 0.21851 dvt2 = 0.04 dvt0w = 7.7
+ dvt1w = 1.272E6 dvt2w = -0.032 vfbsdoff = 0
+ u0 = 4.34156E-2 lu0 = -8.421109E-10 ua = 7.566513E-10
+ lua = 1.068047E-16 ub = 4.96249E-20 lub = -2.461234E-25
+ uc = 3.2583E-11 ud = 0 up = 0
+ lp = 1 eu = 1.67 vsat = 6.660431E4
+ lvsat = 4.347646E-3 a0 = 0.091972 la0 = -1.031265E-8
+ ags = 0.88029 b0 = 3.3993E-7 b1 = 0
+ keta = -0.019904 a1 = 0 a2 = 0.962934
+ rdsw = 430 rdswmin = 0 rdw = 0
+ rdwmin = 0 rsw = 0 rswmin = 0
+ prwb = 0 prwg = 1E-12 wr = 1
+ voff = 0 voffl = 1.944533E-8 minv = 0
+ nfactor = 0.690724 lnfactor = -8.801759E-8 eta0 = 9
+ etab = -2.1692E-4 dsub = 0.42 cit = 9.258412E-8
+ cdsc = 0 cdscb = 1.415095E-7 cdscd = 1.5E-5
+ pclm = 0.11748 pdiblc1 = 8.833E-7 pdiblc2 = 2E-4
+ pdiblcb = 0 drout = 0.13139 pscbe1 = 2.4476E8
+ pscbe2 = 3.84E-9 pvag = 4.541944 delta = 7E-3
+ fprout = 0 pdits = 3.70557E-2 lpdits = -3.174752E-8
+ pditsl = 0 pditsd = 0 lambda = 0
+ vtl = 0 lc = 5E-9 xn = 3
+ alpha0 = 1.950984E-6 lalpha0 = 1.351675E-13 alpha1 = 6.81621E-2
+ lalpha1 = 4.740963E-8 beta0 = 19.026525 lbeta0 = 5.720967E-6
+ aigbacc = 1 bigbacc = 0 cigbacc = 0
+ nigbacc = 1 aigbinv = 0.35 bigbinv = 0.03
+ cigbinv = 6E-3 eigbinv = 1.1 nigbinv = 3
+ aigc = 0.43 bigc = 0.054 cigc = 0.075
+ aigsd = 0.43 bigsd = 0.054 cigsd = 0.075
+ dlcig = 0 nigc = 1 poxedge = 1
+ pigcd = 1 ntox = 1 toxref = 1.16E-8
+ agidl = 0 bgidl = 2.3E9 cgidl = 0.5
+ egidl = 0.8 noia = 2.5E41 noib = 0
+ noic = 0 em = 4.1E7 af = 1
+ ef = 1 kf = 0 lintnoi = 0
+ tnoia = 7.6E6 tnoib = 7.2E6 ntnoi = 1
+ rnoia = 0.8 rnoib = 0.38 xpart = 0
+ cgso = {2.678273E-10/sw_func_tox_hv_ratio} cgdo = {2.678273E-10/sw_func_tox_hv_ratio} cgbo = {0/sw_func_tox_hv_ratio}
+ ckappas = 0.6 cf = 0 clc = 1E-7
+ cle = 0.6 dlc = 6.0712E-8 dwc = 0
+ vfbcv = -1 noff = 4 voffcv = 0.216
+ acde = 1.16 moin = 15 cgsl = {3.85585E-11/sw_func_tox_hv_ratio}
+ cgdl = {3.85585E-11/sw_func_tox_hv_ratio} ijthsrev = 0.1 ijthsfwd = 0.1
+ xjbvs = 1 bvs = 12.69 jss = 4.2966E-4
+ jsws = 8.04E-10 cjs = {8.310E-04*sw_func_nsd_pw_cj} mjs = 0.28329
+ mjsws = 0.057926 cjsws = {8.887314E-11*sw_func_nsd_pw_cj} cjswgs = {3.736446E-11*sw_func_nsd_pw_cj}
+ mjswgs = 0.33 pbs = 0.66345 pbsws = 1
+ pbswgs = 0.2442 xrcrg1 = 12 xrcrg2 = 1
+ rbpb = 50 rbpd = 50 rbps = 50
+ rbdb = 50 rbsb = 50 gbmin = 1E-12
+ tnom = 30 ute = -2.063557 lute = 5.164583E-7
+ kt1 = -0.345969 lkt1 = -2.347392E-8 kt1l = 0
+ kt2 = -1.99578E-2 lkt2 = 7.337204E-9 ua1 = -4.2384E-11
+ lua1 = 8.979096E-16 ub1 = -2.039606E-18 lub1 = 1.142911E-24
+ uc1 = -8.195316E-11 luc1 = 7.920845E-17 at = 4.805277E3
+ lat = 1.26477E-2 prt = 0 njs = 1.5764
+ xtis = 0 tpb = 1.9685E-3 tpbsw = 1E-3
+ tpbswg = 0 tcj = 8.3E-4 tcjsw = 0
+ tcjswg = 0 tvoff = 0 tvfbsdoff = 0
+ saref = 3E-6 sbref = 3E-6 wlod = 0
+ ku0 = -3E-8 kvsat = 0.4 kvth0 = -7E-9
+ tku0 = 0 llodku0 = 0 wlodku0 = 1
+ llodvth = 0 wlodvth = 1 lku0 = 0
+ wku0 = 2E-7 pku0 = 0 lkvth0 = 0
+ wkvth0 = 8E-7 pkvth0 = 0 stk2 = 0
+ lodk2 = 1 steta0 = 0 lodeta0 = 1

.model nhvnative_model.5 nmos
+ level = 54 lmin = 9E-7 lmax = 1E-6 wmin = 1E-5
+ wmax = 1.01E-4 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 1.16E-8
+ toxm = 1.16E-8 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 1E23 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {4.5E-8+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {6.93E-8-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = -4.6E-9 dwb = 1.92E-9 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = 6.08069E-2 k1 = 0.364
+ k2 = 4.04085E-2 k3 = 1.4 k3b = -0.58
+ w0 = 0 lpe0 = -1.236227E-14 lpeb = 0
+ vbm = -3 dvtp0 = 0 dvtp1 = 0
+ dvt0 = 5.7 dvt1 = 0.21851 dvt2 = 0.04
+ dvt0w = 7.7 dvt1w = 1.272E6 dvt2w = -0.032
+ vfbsdoff = 0 u0 = 0.042438 ua = 8.80641E-10
+ ub = -2.361E-19 uc = 3.2583E-11 ud = 0
+ up = 0 lp = 1 eu = 1.67
+ vsat = 7.16515E4 a0 = 0.08 ags = 0.87995
+ b0 = 3.3993E-7 b1 = 0 keta = -0.019904
+ a1 = 0 a2 = 0.962934 rdsw = 430
+ rdswmin = 0 rdw = 0 rdwmin = 0
+ rsw = 0 rswmin = 0 prwb = 0
+ prwg = 1E-12 wr = 1 voff = 0
+ voffl = 1.944533E-8 minv = 0 nfactor = 0.588544
+ eta0 = 9 etab = -2.1692E-4 dsub = 0.42
+ cit = 9.258412E-8 cdsc = 0 cdscb = 1.415095E-7
+ cdscd = 1.5E-5 pclm = 0.11748 pdiblc1 = 8.833E-7
+ pdiblc2 = 2E-4 pdiblcb = 0 drout = 0.13139
+ pscbe1 = 2.4476E8 pscbe2 = 3.84E-9 pvag = 4.541944
+ delta = 7E-3 fprout = 0 pdits = 2E-4
+ pditsl = 0 pditsd = 0 lambda = 0
+ vtl = 0 lc = 5E-9 xn = 3
+ alpha0 = 2.1079E-6 alpha1 = 0.1232 beta0 = 25.668
+ aigbacc = 1 bigbacc = 0 cigbacc = 0
+ nigbacc = 1 aigbinv = 0.35 bigbinv = 0.03
+ cigbinv = 6E-3 eigbinv = 1.1 nigbinv = 3
+ aigc = 0.43 bigc = 0.054 cigc = 0.075
+ aigsd = 0.43 bigsd = 0.054 cigsd = 0.075
+ dlcig = 0 nigc = 1 poxedge = 1
+ pigcd = 1 ntox = 1 toxref = 1.16E-8
+ agidl = 0 bgidl = 2.3E9 cgidl = 0.5
+ egidl = 0.8 noia = 2.5E41 noib = 0
+ noic = 0 em = 4.1E7 af = 1
+ ef = 1 kf = 0 lintnoi = 0
+ tnoia = 7.6E6 tnoib = 7.2E6 ntnoi = 1
+ rnoia = 0.8 rnoib = 0.38 xpart = 0
+ cgso = {2.678273E-10/sw_func_tox_hv_ratio} cgdo = {2.678273E-10/sw_func_tox_hv_ratio} cgbo = {0/sw_func_tox_hv_ratio}
+ ckappas = 0.6 cf = 0 clc = 1E-7
+ cle = 0.6 dlc = 6.0712E-8 dwc = 0
+ vfbcv = -1 noff = 4 voffcv = 0.216
+ acde = 1.16 moin = 15 cgsl = {3.85585E-11/sw_func_tox_hv_ratio}
+ cgdl = {3.85585E-11/sw_func_tox_hv_ratio} ijthsrev = 0.1 ijthsfwd = 0.1
+ xjbvs = 1 bvs = 12.69 jss = 4.2966E-4
+ jsws = 8.04E-10 cjs = {8.310E-04*sw_func_nsd_pw_cj} mjs = 0.28329
+ mjsws = 0.057926 cjsws = {8.887314E-11*sw_func_nsd_pw_cj} cjswgs = {3.736446E-11*sw_func_nsd_pw_cj}
+ mjswgs = 0.33 pbs = 0.66345 pbsws = 1
+ pbswgs = 0.2442 xrcrg1 = 12 xrcrg2 = 1
+ rbpb = 50 rbpd = 50 rbps = 50
+ rbdb = 50 rbsb = 50 gbmin = 1E-12
+ tnom = 30 ute = -1.464 kt1 = -0.37322
+ kt1l = 0 kt2 = -0.01144 ua1 = 1E-9
+ ub1 = -7.128E-19 uc1 = 1E-11 at = 1.9488E4
+ prt = 0 njs = 1.5764 xtis = 0
+ tpb = 1.9685E-3 tpbsw = 1E-3 tpbswg = 0
+ tcj = 8.3E-4 tcjsw = 0 tcjswg = 0
+ tvoff = 0 tvfbsdoff = 0 saref = 2.54E-6
+ sbref = 2.54E-6 wlod = 0 ku0 = -3E-8
+ kvsat = 0.4 kvth0 = -7E-9 tku0 = 0
+ llodku0 = 0 wlodku0 = 1 llodvth = 0
+ wlodvth = 1 lku0 = 0 wku0 = 2E-7
+ pku0 = 0 lkvth0 = 0 wkvth0 = 8E-7
+ pkvth0 = 0 stk2 = 0 lodk2 = 1
+ steta0 = 0 lodeta0 = 1

.model nhvnative_model.6 nmos
+ level = 54 lmin = 8E-6 lmax = 2.525E-5 wmin = 1E-6
+ wmax = 1E-5 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 1.16E-8
+ toxm = 1.16E-8 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 1E23 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {4.5E-8+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {6.93E-8-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = -4.6E-9 dwb = 1.92E-9 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = 0.038459 lvth0 = 2.72244E-8
+ k1 = 0.364 k2 = 0.041446 lk2 = -1.271545E-8
+ k3 = 1.4 k3b = -0.58 w0 = 0
+ lpe0 = -1.236227E-14 lpeb = 0 vbm = -3
+ dvtp0 = 0 dvtp1 = 0 dvt0 = 5.7
+ dvt1 = 0.21851 dvt2 = 0.04 dvt0w = 7.7
+ dvt1w = 1.272E6 dvt2w = -0.032 vfbsdoff = 0
+ u0 = 4.45181E-2 lu0 = -2.145301E-9 ua = 1.096856E-9
+ lua = -2.413176E-17 ub = -1.500717E-19 lub = -1.033446E-24
+ uc = 1.9159E-11 ud = 0 up = 0
+ lp = 1 eu = 1.67 vsat = 7.5917E4
+ a0 = 1.387857 la0 = -1.035676E-5 ags = 2.90552E-2
+ lags = 3.780528E-6 b0 = 5.734E-8 b1 = 4.9905E-8
+ keta = -7.522213E-3 lketa = -1.067247E-7 a1 = 0
+ a2 = 0.962934 rdsw = 430 rdswmin = 0
+ rdw = 0 rdwmin = 0 rsw = 0
+ rswmin = 0 prwb = 0 prwg = 1E-12
+ wr = 1 voff = 0 voffl = 1.944533E-8
+ minv = 0 nfactor = 0.701166 lnfactor = -9.975764E-8
+ eta0 = 9 etab = -2.1692E-4 dsub = 0.42
+ cit = 9.258412E-8 cdsc = 0 cdscb = 1.415095E-7
+ cdscd = 1.5E-5 pclm = 0.089 pdiblc1 = 1.0772E-6
+ pdiblc2 = 5.1E-4 pdiblcb = 0 drout = 0.11135
+ pscbe1 = 2.7814E8 pscbe2 = 1.6E-8 pvag = 4.541944
+ delta = 7E-3 fprout = 0 pdits = -2.630332E-3
+ lpdits = 6.539373E-8 pditsl = 0 pditsd = 0
+ lambda = 0 vtl = 0 lc = 5E-9
+ xn = 3 alpha0 = 2.97923E-6 lalpha0 = -2.08346E-11
+ alpha1 = 0.5456 beta0 = 20.117451 lbeta0 = -8.73756E-6
+ aigbacc = 1 bigbacc = 0 cigbacc = 0
+ nigbacc = 1 aigbinv = 0.35 bigbinv = 0.03
+ cigbinv = 6E-3 eigbinv = 1.1 nigbinv = 3
+ aigc = 0.43 bigc = 0.054 cigc = 0.075
+ aigsd = 0.43 bigsd = 0.054 cigsd = 0.075
+ dlcig = 0 nigc = 1 poxedge = 1
+ pigcd = 1 ntox = 1 toxref = 1.16E-8
+ agidl = 0 bgidl = 2.3E9 cgidl = 0.5
+ egidl = 0.8 noia = 2.5E41 noib = 0
+ noic = 0 em = 4.1E7 af = 1
+ ef = 1 kf = 0 lintnoi = 0
+ tnoia = 7.6E6 tnoib = 7.2E6 ntnoi = 1
+ rnoia = 0.8 rnoib = 0.38 xpart = 0
+ cgso = {2.678273E-10/sw_func_tox_hv_ratio} cgdo = {2.678273E-10/sw_func_tox_hv_ratio} cgbo = {0/sw_func_tox_hv_ratio}
+ ckappas = 0.6 cf = 0 clc = 1E-7
+ cle = 0.6 dlc = 6.0712E-8 dwc = 0
+ vfbcv = -1 noff = 4 voffcv = 0.216
+ acde = 1.16 moin = 15 cgsl = {3.85585E-11/sw_func_tox_hv_ratio}
+ cgdl = {3.85585E-11/sw_func_tox_hv_ratio} ijthsrev = 0.1 ijthsfwd = 0.1
+ xjbvs = 1 bvs = 12.69 jss = 4.2966E-4
+ jsws = 8.04E-10 cjs = {8.310E-04*sw_func_nsd_pw_cj} mjs = 0.28329
+ mjsws = 0.057926 cjsws = {8.887314E-11*sw_func_nsd_pw_cj} cjswgs = {3.736446E-11*sw_func_nsd_pw_cj}
+ mjswgs = 0.33 pbs = 0.66345 pbsws = 1
+ pbswgs = 0.2442 xrcrg1 = 12 xrcrg2 = 1
+ rbpb = 50 rbpd = 50 rbps = 50
+ rbdb = 50 rbsb = 50 gbmin = 1E-12
+ tnom = 30 ute = -1.464 kt1 = -0.370524
+ lkt1 = 1.149679E-7 kt1l = 0 kt2 = -0.01144
+ ua1 = 1E-9 ub1 = -1.088076E-18 lub1 = 2.950191E-24
+ uc1 = 1E-11 at = 8.63772E4 lat = -0.496661
+ prt = 0 njs = 1.5764 xtis = 0
+ tpb = 1.9685E-3 tpbsw = 1E-3 tpbswg = 0
+ tcj = 8.3E-4 tcjsw = 0 tcjswg = 0
+ tvoff = 0 tvfbsdoff = 0 saref = 3E-6
+ sbref = 3E-6 wlod = 0 ku0 = -3E-8
+ kvsat = 0.4 kvth0 = -7E-9 tku0 = 0
+ llodku0 = 0 wlodku0 = 1 llodvth = 0
+ wlodvth = 1 lku0 = 0 wku0 = 2E-7
+ pku0 = 0 lkvth0 = 0 wkvth0 = 8E-7
+ pkvth0 = 0 stk2 = 0 lodk2 = 1
+ steta0 = 0 lodeta0 = 1

.model nhvnative_model.7 nmos
+ level = 54 lmin = 4E-6 lmax = 8E-6 wmin = 1E-6
+ wmax = 1E-5 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 1.16E-8
+ toxm = 1.16E-8 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 1E23 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {4.5E-8+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {6.93E-8-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = -4.6E-9 dwb = 1.92E-9 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = 2.46565E-2 lvth0 = 1.357307E-7
+ wvth0 = 1.920393E-8 pvth0 = -1.509698E-13 k1 = 0.364
+ k2 = 4.00866E-2 lk2 = -2.029296E-9 wk2 = 5.548674E-10
+ pk2 = -4.362034E-15 k3 = 1.4 k3b = -0.58
+ w0 = 0 lpe0 = -1.236227E-14 lpeb = 0
+ vbm = -3 dvtp0 = 0 dvtp1 = 0
+ dvt0 = 5.7 dvt1 = 0.21851 dvt2 = 0.04
+ dvt0w = 7.7 dvt1w = 1.272E6 dvt2w = -0.032
+ vfbsdoff = 0 u0 = 0.045857 lu0 = -1.267135E-8
+ wu0 = -1.435944E-9 pu0 = 1.128853E-14 ua = 1.388192E-9
+ lua = -2.314443E-15 wua = -2.657246E-16 pua = 2.088968E-21
+ ub = -5.714349E-19 lub = 2.279058E-24 wub = 2.982933E-25
+ pub = -2.345003E-30 uc = 6.745028E-12 luc = 9.75912E-17
+ wuc = 1.954035E-17 puc = -1.536145E-22 ud = 0
+ up = 0 lp = 1 eu = 1.67
+ vsat = 7.879152E4 lvsat = -2.25978E-2 wvsat = -1.307778E-3
+ pvsat = 1.028097E-8 a0 = 5.99938E-2 la0 = 8.209869E-8
+ wa0 = -1.437601E-8 pa0 = 1.130156E-13 ags = 0.304895
+ lags = 1.612045E-6 wags = 1.815598E-7 pags = -1.427315E-12
+ b0 = -2.576375E-7 lb0 = 2.476164E-12 wb0 = 4.179966E-13
+ pb0 = -3.286039E-18 b1 = 1.029519E-7 lb1 = -4.170229E-13
+ wb1 = -4.827268E-14 pb1 = 3.794908E-19 keta = -2.23672E-2
+ lketa = 9.977464E-9 wketa = 1.154946E-9 pketa = -9.079492E-15
+ a1 = 0 a2 = 0.962934 rdsw = 430
+ rdswmin = 0 rdw = 0 rdwmin = 0
+ rsw = 0 rswmin = 0 prwb = 0
+ prwg = 1E-12 wr = 1 voff = 0
+ voffl = 1.944533E-8 minv = 0 nfactor = 0.715248
+ lnfactor = -2.104628E-7 wnfactor = -2.237248E-8 pnfactor = 1.75879E-13
+ eta0 = 9 etab = -2.1692E-4 dsub = 0.42
+ cit = 9.258412E-8 cdsc = 0 cdscb = 1.415095E-7
+ cdscd = 1.5E-5 pclm = 0.058727 lpclm = 2.379884E-7
+ wpclm = 2.754846E-8 ppclm = -2.165695E-13 pdiblc1 = 1.283307E-6
+ lpdiblc1 = -1.620293E-12 wpdiblc1 = -1.875578E-13 ppdiblc1 = 1.474467E-18
+ pdiblc2 = 8.395169E-4 lpdiblc2 = -2.590464E-9 wpdiblc2 = -2.998603E-10
+ ppdiblc2 = 2.357322E-15 pdiblcb = 0 drout = 9.00483E-2
+ ldrout = 1.67461E-7 wdrout = 1.938452E-8 pdrout = -1.523895E-13
+ pscbe1 = 3.136215E8 lpscbe1 = -278.934461 wpscbe1 = -32.288188
+ ppscbe1 = 2.538304E-4 pscbe2 = 2.892556E-8 lpscbe2 = -1.01613E-13
+ wpscbe2 = -1.176226E-14 ppscbe2 = 9.246786E-20 pvag = 4.541944
+ delta = 7E-3 fprout = 0 pdits = 4.505991E-3
+ lpdits = 9.292244E-9 wpdits = 1.075628E-9 ppdits = -8.455942E-15
+ pditsl = 0 pditsd = 0 lambda = 0
+ vtl = 0 lc = 5E-9 xn = 3
+ alpha0 = -1.457852E-6 lalpha0 = 1.404708E-11 walpha0 = 1.626027E-12
+ palpha0 = -1.278285E-17 alpha1 = 1.026023 lalpha1 = -3.776796E-6
+ walpha1 = -4.371848E-7 palpha1 = 3.436884E-12 beta0 = 18.536173
+ lbeta0 = 3.6935E-6 wbeta0 = 4.275428E-7 pbeta0 = -3.361085E-12
+ aigbacc = 1 bigbacc = 0 cigbacc = 0
+ nigbacc = 1 aigbinv = 0.35 bigbinv = 0.03
+ cigbinv = 6E-3 eigbinv = 1.1 nigbinv = 3
+ aigc = 0.43 bigc = 0.054 cigc = 0.075
+ aigsd = 0.43 bigsd = 0.054 cigsd = 0.075
+ dlcig = 0 nigc = 1 poxedge = 1
+ pigcd = 1 ntox = 1 toxref = 1.16E-8
+ agidl = 0 bgidl = 2.3E9 cgidl = 0.5
+ egidl = 0.8 noia = 2.5E41 noib = 0
+ noic = 0 em = 4.1E7 af = 1
+ ef = 1 kf = 0 lintnoi = 0
+ tnoia = 7.6E6 tnoib = 7.2E6 ntnoi = 1
+ rnoia = 0.8 rnoib = 0.38 xpart = 0
+ cgso = {2.678273E-10/sw_func_tox_hv_ratio} cgdo = {2.678273E-10/sw_func_tox_hv_ratio} cgbo = {0/sw_func_tox_hv_ratio}
+ ckappas = 0.6 cf = 0 clc = 1E-7
+ cle = 0.6 dlc = 6.0712E-8 dwc = 0
+ vfbcv = -1 noff = 4 voffcv = 0.216
+ acde = 1.16 moin = 15 cgsl = {3.85585E-11/sw_func_tox_hv_ratio}
+ cgdl = {3.85585E-11/sw_func_tox_hv_ratio} ijthsrev = 0.1 ijthsfwd = 0.1
+ xjbvs = 1 bvs = 12.69 jss = 4.2966E-4
+ jsws = 8.04E-10 cjs = {8.310E-04*sw_func_nsd_pw_cj} mjs = 0.28329
+ mjsws = 0.057926 cjsws = {8.887314E-11*sw_func_nsd_pw_cj} cjswgs = {3.736446E-11*sw_func_nsd_pw_cj}
+ mjswgs = 0.33 pbs = 0.66345 pbsws = 1
+ pbswgs = 0.2442 xrcrg1 = 12 xrcrg2 = 1
+ rbpb = 50 rbpd = 50 rbps = 50
+ rbdb = 50 rbsb = 50 gbmin = 1E-12
+ tnom = 30 ute = -1.121621 lute = -2.691575E-6
+ wute = -3.115646E-7 pute = 2.449334E-12 kt1 = -0.352949
+ lkt1 = -2.320068E-8 wkt1 = -3.607997E-9 pkt1 = 2.836391E-14
+ kt1l = 0 kt2 = -6.575906E-3 lkt2 = -3.823859E-8
+ wkt2 = -4.426326E-9 pkt2 = 3.479712E-14 ua1 = 1.595256E-9
+ lua1 = -4.679548E-15 wua1 = -5.416832E-16 pua1 = 4.258388E-21
+ ub1 = 2.570425E-19 lub1 = -7.62432E-24 wub1 = -8.825567E-25
+ pub1 = 6.938131E-30 uc1 = 6.251011E-11 luc1 = -4.128029E-16
+ wuc1 = -4.77842E-17 puc1 = 3.756507E-22 at = 2.362518E4
+ lat = -3.342534E-3 wat = -3.869166E-4 pat = 3.041706E-9
+ prt = 0 njs = 1.5764 xtis = 0
+ tpb = 1.9685E-3 tpbsw = 1E-3 tpbswg = 0
+ tcj = 8.3E-4 tcjsw = 0 tcjswg = 0
+ tvoff = 0 tvfbsdoff = 0 saref = 3E-6
+ sbref = 3E-6 wlod = 0 ku0 = -3E-8
+ kvsat = 0.4 kvth0 = -7E-9 tku0 = 0
+ llodku0 = 0 wlodku0 = 1 llodvth = 0
+ wlodvth = 1 lku0 = 0 wku0 = 2E-7
+ pku0 = 0 lkvth0 = 0 wkvth0 = 8E-7
+ pkvth0 = 0 stk2 = 0 lodk2 = 1
+ steta0 = 0 lodeta0 = 1

.model nhvnative_model.8 nmos
+ level = 54 lmin = 2E-6 lmax = 4E-6 wmin = 1E-6
+ wmax = 1E-5 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 1.16E-8
+ toxm = 1.16E-8 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 1E23 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {4.5E-8+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {6.93E-8-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = -4.6E-9 dwb = 1.92E-9 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = 6.85342E-2 lvth0 = -3.369843E-8
+ wvth0 = -1.965076E-8 pvth0 = -9.362685E-16 k1 = 0.364
+ k2 = 4.03815E-2 lk2 = -3.167733E-9 wk2 = -5.364654E-12
+ pk2 = -2.198754E-15 k3 = 1.4 k3b = -0.58
+ w0 = 0 lpe0 = -1.236227E-14 lpeb = 0
+ vbm = -3 dvtp0 = 0 dvtp1 = 0
+ dvt0 = 5.7 dvt1 = 0.21851 dvt2 = 0.04
+ dvt0w = 7.7 dvt1w = 1.272E6 dvt2w = -0.032
+ vfbsdoff = 0 u0 = 4.23408E-2 lu0 = 9.063956E-10
+ wu0 = 1.622242E-9 pu0 = -5.203492E-16 ua = 7.911728E-10
+ lua = -9.112971E-18 wua = 2.75477E-16 pua = -8.282375E-25
+ ub = 7.94614E-20 lub = -2.343127E-25 wub = -2.628752E-25
+ pub = -1.781071E-31 uc = 2.934689E-11 luc = 1.031636E-17
+ wuc = -1.781051E-17 puc = -9.387892E-24 ud = 0
+ up = 0 lp = 1 eu = 1.67
+ vsat = 7.778693E4 lvsat = -1.87186E-2 wvsat = -8.538002E-3
+ pvsat = 3.819975E-8 a0 = 7.15327E-2 la0 = 3.754209E-8
+ wa0 = 7.735645E-8 pa0 = -2.412001E-13 ags = 0.539788
+ lags = 7.050256E-7 wags = -1.024506E-8 pags = -6.866791E-13
+ b0 = 3.836232E-7 wb0 = -4.330001E-13 b1 = -5.04595E-9
+ wb1 = 5.000536E-14 keta = -1.97833E-2 wketa = -1.196401E-9
+ a1 = 0 a2 = 0.962934 rdsw = 430
+ rdswmin = 0 rdw = 0 rdwmin = 0
+ rsw = 0 rswmin = 0 prwb = 0
+ prwg = 1E-12 wr = 1 voff = 0
+ voffl = 1.944533E-8 minv = 0 nfactor = 0.678175
+ lnfactor = -6.731035E-8 wnfactor = 3.160969E-8 pnfactor = -3.256774E-14
+ eta0 = 9 etab = -2.1692E-4 dsub = 0.42
+ cit = 9.258412E-8 cdsc = 0 cdscb = 1.415095E-7
+ cdscd = 1.5E-5 pclm = 0.12036 wpclm = -2.853728E-8
+ pdiblc1 = 8.636946E-7 wpdiblc1 = 1.9429E-13 pdiblc2 = 1.686556E-4
+ wpdiblc2 = 3.106234E-10 pdiblcb = 0 drout = 0.133416
+ wdrout = -2.00803E-8 pscbe1 = 2.413849E8 wpscbe1 = 33.447131
+ pscbe2 = 2.610489E-9 wpscbe2 = 1.218446E-14 pvag = 4.541944
+ delta = 7E-3 fprout = 0 pdits = -5.663398E-3
+ lpdits = 4.856032E-8 wpdits = 1.765545E-9 ppdits = -1.111999E-14
+ pditsl = 0 pditsd = 0 lambda = 0
+ vtl = 0 lc = 5E-9 xn = 3
+ alpha0 = 2.307066E-6 lalpha0 = -4.90774E-13 walpha0 = -3.069362E-12
+ palpha0 = 5.347929E-18 alpha1 = 0.047933 walpha1 = 4.52877E-7
+ beta0 = 17.066069 lbeta0 = 9.37016E-6 wbeta0 = -8.550856E-7
+ pbeta0 = 1.591656E-12 aigbacc = 1 bigbacc = 0
+ cigbacc = 0 nigbacc = 1 aigbinv = 0.35
+ bigbinv = 0.03 cigbinv = 6E-3 eigbinv = 1.1
+ nigbinv = 3 aigc = 0.43 bigc = 0.054
+ cigc = 0.075 aigsd = 0.43 bigsd = 0.054
+ cigsd = 0.075 dlcig = 0 nigc = 1
+ poxedge = 1 pigcd = 1 ntox = 1
+ toxref = 1.16E-8 agidl = 0 bgidl = 2.3E9
+ cgidl = 0.5 egidl = 0.8 noia = 2.5E41
+ noib = 0 noic = 0 em = 4.1E7
+ af = 1 ef = 1 kf = 0
+ lintnoi = 0 tnoia = 7.6E6 tnoib = 7.2E6
+ ntnoi = 1 rnoia = 0.8 rnoib = 0.38
+ xpart = 0 cgso = {2.678273E-10/sw_func_tox_hv_ratio} cgdo = {2.678273E-10/sw_func_tox_hv_ratio}
+ cgbo = {0/sw_func_tox_hv_ratio} ckappas = 0.6 cf = 0
+ clc = 1E-7 cle = 0.6 dlc = 6.0712E-8
+ dwc = 0 vfbcv = -1 noff = 4
+ voffcv = 0.216 acde = 1.16 moin = 15
+ cgsl = {3.85585E-11/sw_func_tox_hv_ratio} cgdl = {3.85585E-11/sw_func_tox_hv_ratio} ijthsrev = 0.1
+ ijthsfwd = 0.1 xjbvs = 1 bvs = 12.69
+ jss = 4.2966E-4 jsws = 8.04E-10 cjs = {8.310E-04*sw_func_nsd_pw_cj}
+ mjs = 0.28329 mjsws = 0.057926 cjsws = {8.887314E-11*sw_func_nsd_pw_cj}
+ cjswgs = {3.736446E-11*sw_func_nsd_pw_cj} mjswgs = 0.33 pbs = 0.66345
+ pbsws = 1 pbswgs = 0.2442 xrcrg1 = 12
+ xrcrg2 = 1 rbpb = 50 rbpd = 50
+ rbps = 50 rbdb = 50 rbsb = 50
+ gbmin = 1E-12 tnom = 30 ute = -1.818668
+ wute = 3.227478E-7 kt1 = -0.359997 lkt1 = 4.015278E-9
+ wkt1 = 1.404242E-8 pkt1 = -3.979141E-14 kt1l = 0
+ kt2 = -1.64787E-2 wkt2 = 4.585203E-9 ua1 = 3.833778E-10
+ wua1 = 5.611262E-16 ub1 = -1.922005E-18 lub1 = 7.898528E-25
+ wub1 = 1.100376E-24 pub1 = -7.187661E-31 uc1 = -4.439489E-11
+ wuc1 = 4.949935E-17 at = 3.29711E4 lat = -3.94308E-2
+ wat = 2.504686E-3 pat = -8.123929E-9 prt = 0
+ njs = 1.5764 xtis = 0 tpb = 1.9685E-3
+ tpbsw = 1E-3 tpbswg = 0 tcj = 8.3E-4
+ tcjsw = 0 tcjswg = 0 tvoff = 0
+ tvfbsdoff = 0 saref = 3E-6 sbref = 3E-6
+ wlod = 0 ku0 = -3E-8 kvsat = 0.4
+ kvth0 = -7E-9 tku0 = 0 llodku0 = 0
+ wlodku0 = 1 llodvth = 0 wlodvth = 1
+ lku0 = 0 wku0 = 2E-7 pku0 = 0
+ lkvth0 = 0 wkvth0 = 8E-7 pkvth0 = 0
+ stk2 = 0 lodk2 = 1 steta0 = 0
+ lodeta0 = 1

.model nhvnative_model.9 nmos
+ level = 54 lmin = 1E-6 lmax = 2E-6 wmin = 1E-6
+ wmax = 1E-5 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 1.16E-8
+ toxm = 1.16E-8 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 1E23 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {4.5E-8+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {6.93E-8-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = -4.6E-9 dwb = 1.92E-9 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = 3.94835E-2 lvth0 = 2.037651E-8
+ wvth0 = -1.760958E-8 pvth0 = -4.735716E-15 k1 = 0.364
+ k2 = 3.71041E-2 lk2 = 2.932735E-9 wk2 = -1.353221E-9
+ pk2 = 3.101447E-16 k3 = 1.4 k3b = -0.58
+ w0 = 0 lpe0 = -1.236227E-14 lpeb = 0
+ vbm = -3 dvtp0 = 0 dvtp1 = 0
+ dvt0 = 5.7 dvt1 = 0.21851 dvt2 = 0.04
+ dvt0w = 7.7 dvt1w = 1.272E6 dvt2w = -0.032
+ vfbsdoff = 0 u0 = 4.32808E-2 lu0 = -8.434565E-10
+ wu0 = 1.335531E-9 pu0 = 1.333507E-17 ua = 7.226882E-10
+ lua = 1.183642E-16 wua = 3.365742E-16 pua = -1.145547E-22
+ ub = 8.701715E-20 lub = -2.483769E-25 wub = -3.705572E-25
+ pub = 2.233222E-32 uc = 3.488915E-11 wuc = -2.285397E-17
+ ud = 0 up = 0 lp = 1
+ eu = 1.67 vsat = 6.523529E4 lvsat = 4.644979E-3
+ wvsat = 0.013567 pvsat = -2.946568E-9 a0 = 0.10091
+ la0 = -1.714104E-8 wa0 = -8.857753E-8 pa0 = 6.766936E-14
+ ags = 0.91961 lags = -1.973462E-9 wags = -3.867528E-7
+ pags = 1.415241E-14 b0 = 3.836232E-7 wb0 = -4.330001E-13
+ b1 = -5.04595E-9 wb1 = 5.000536E-14 keta = -1.97833E-2
+ wketa = -1.196401E-9 a1 = 0 a2 = 0.962934
+ rdsw = 430 rdswmin = 0 rdw = 0
+ rdwmin = 0 rsw = 0 rswmin = 0
+ prwb = 0 prwg = 1E-12 wr = 1
+ voff = 0 voffl = 1.944533E-8 minv = 0
+ nfactor = 0.692098 lnfactor = -9.322623E-8 wnfactor = -1.361722E-8
+ pnfactor = 5.161763E-14 eta0 = 9 etab = -2.1692E-4
+ dsub = 0.42 cit = 9.258412E-8 cdsc = 0
+ cdscb = 1.415095E-7 cdscd = 1.5E-5 pclm = 0.12036
+ wpclm = -2.853728E-8 pdiblc1 = 8.636946E-7 wpdiblc1 = 1.9429E-13
+ pdiblc2 = 1.24236E-4 lpdiblc2 = 8.268251E-11 wpdiblc2 = 7.50821E-10
+ ppdiblc2 = -8.193836E-16 pdiblcb = 0 drout = 0.133416
+ wdrout = -2.00803E-8 pscbe1 = 2.413849E8 wpscbe1 = 33.447131
+ pscbe2 = 2.610489E-9 wpscbe2 = 1.218446E-14 pvag = 4.541944
+ delta = 7E-3 fprout = 0 pdits = 3.78288E-2
+ lpdits = -3.239601E-8 wpdits = -7.660976E-9 ppdits = 6.426538E-15
+ pditsl = 0 pditsd = 0 lambda = 0
+ vtl = 0 lc = 5E-9 xn = 3
+ alpha0 = 1.963449E-6 lalpha0 = 1.488344E-13 walpha0 = -1.235319E-13
+ palpha0 = -1.354393E-19 alpha1 = 1.98879E-2 lalpha1 = 5.220327E-8
+ walpha1 = 4.783981E-7 palpha1 = -4.750497E-14 beta0 = 18.930892
+ lbeta0 = 5.898977E-6 wbeta0 = 9.477193E-7 pbeta0 = -1.764085E-12
+ aigbacc = 1 bigbacc = 0 cigbacc = 0
+ nigbacc = 1 aigbinv = 0.35 bigbinv = 0.03
+ cigbinv = 6E-3 eigbinv = 1.1 nigbinv = 3
+ aigc = 0.43 bigc = 0.054 cigc = 0.075
+ aigsd = 0.43 bigsd = 0.054 cigsd = 0.075
+ dlcig = 0 nigc = 1 poxedge = 1
+ pigcd = 1 ntox = 1 toxref = 1.16E-8
+ agidl = 0 bgidl = 2.3E9 cgidl = 0.5
+ egidl = 0.8 noia = 2.5E41 noib = 0
+ noic = 0 em = 4.1E7 af = 1
+ ef = 1 kf = 0 lintnoi = 0
+ tnoia = 7.6E6 tnoib = 7.2E6 ntnoi = 1
+ rnoia = 0.8 rnoib = 0.38 xpart = 0
+ cgso = {2.678273E-10/sw_func_tox_hv_ratio} cgdo = {2.678273E-10/sw_func_tox_hv_ratio} cgbo = {0/sw_func_tox_hv_ratio}
+ ckappas = 0.6 cf = 0 clc = 1E-7
+ cle = 0.6 dlc = 6.0712E-8 dwc = 0
+ vfbcv = -1 noff = 4 voffcv = 0.216
+ acde = 1.16 moin = 15 cgsl = {3.85585E-11/sw_func_tox_hv_ratio}
+ cgdl = {3.85585E-11/sw_func_tox_hv_ratio} ijthsrev = 0.1 ijthsfwd = 0.1
+ xjbvs = 1 bvs = 12.69 jss = 4.2966E-4
+ jsws = 8.04E-10 cjs = {8.310E-04*sw_func_nsd_pw_cj} mjs = 0.28329
+ mjsws = 0.057926 cjsws = {8.887314E-11*sw_func_nsd_pw_cj} cjswgs = {3.736446E-11*sw_func_nsd_pw_cj}
+ mjswgs = 0.33 pbs = 0.66345 pbsws = 1
+ pbswgs = 0.2442 xrcrg1 = 12 xrcrg2 = 1
+ rbpb = 50 rbpd = 50 rbps = 50
+ rbdb = 50 rbsb = 50 gbmin = 1E-12
+ tnom = 30 ute = -2.124179 lute = 5.68678E-7
+ wute = 6.007627E-7 pute = -5.17497E-13 kt1 = -0.343954
+ lkt1 = -2.58474E-8 wkt1 = -1.997098E-8 pkt1 = 2.352113E-14
+ kt1l = 0 kt2 = -0.020819 lkt2 = 8.079077E-9
+ wkt2 = 8.534897E-9 pkt2 = -7.35196E-15 ua1 = -1.477806E-10
+ lua1 = 9.886982E-16 wua1 = 1.04448E-15 pua1 = -8.997154E-22
+ ub1 = -2.173761E-18 lub1 = 1.258472E-24 wub1 = 1.329474E-24
+ pub1 = -1.145209E-30 uc1 = -9.125065E-11 luc1 = 8.721731E-17
+ wuc1 = 9.213809E-17 puc1 = -7.936775E-23 at = 5.195004E3
+ lat = 1.22716E-2 wat = -3.8622E-3 pat = 3.727392E-9
+ prt = 0 njs = 1.5764 xtis = 0
+ tpb = 1.9685E-3 tpbsw = 1E-3 tpbswg = 0
+ tcj = 8.3E-4 tcjsw = 0 tcjswg = 0
+ tvoff = 0 tvfbsdoff = 0 saref = 3E-6
+ sbref = 3E-6 wlod = 0 ku0 = -3E-8
+ kvsat = 0.4 kvth0 = -7E-9 tku0 = 0
+ llodku0 = 0 wlodku0 = 1 llodvth = 0
+ wlodvth = 1 lku0 = 0 wku0 = 2E-7
+ pku0 = 0 lkvth0 = 0 wkvth0 = 8E-7
+ pkvth0 = 0 stk2 = 0 lodk2 = 1
+ steta0 = 0 lodeta0 = 1

.model nhvnative_model.10 nmos
+ level = 54 lmin = 9E-7 lmax = 1E-6 wmin = 1E-6
+ wmax = 1E-5 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 1.16E-8
+ toxm = 1.16E-8 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 1E23 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {4.5E-8+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {6.93E-8-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = -4.6E-9 dwb = 1.92E-9 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = 6.31386E-2 wvth0 = -2.310728E-8
+ k1 = 0.364 k2 = 4.05087E-2 wk2 = -9.931734E-10
+ k3 = 1.4 k3b = -0.58 w0 = 0
+ lpe0 = -1.236227E-14 lpeb = 0 vbm = -3
+ dvtp0 = 0 dvtp1 = 0 dvt0 = 5.7
+ dvt1 = 0.21851 dvt2 = 0.04 dvt0w = 7.7
+ dvt1w = 1.272E6 dvt2w = -0.032 vfbsdoff = 0
+ u0 = 4.23017E-2 wu0 = 1.351012E-9 ua = 8.600973E-10
+ wua = 2.035876E-16 ub = -2.013238E-19 wub = -3.446317E-25
+ uc = 3.488915E-11 wuc = -2.285397E-17 ud = 0
+ up = 0 lp = 1 eu = 1.67
+ vsat = 7.062765E4 wvsat = 1.01464E-2 a0 = 8.10111E-2
+ wa0 = -1.002011E-8 ags = 0.917319 wags = -3.703233E-7
+ b0 = 3.836232E-7 wb0 = -4.330001E-13 b1 = -5.04595E-9
+ wb1 = 5.000536E-14 keta = -1.97833E-2 wketa = -1.196401E-9
+ a1 = 0 a2 = 0.962934 rdsw = 430
+ rdswmin = 0 rdw = 0 rdwmin = 0
+ rsw = 0 rswmin = 0 prwb = 0
+ prwg = 1E-12 wr = 1 voff = 0
+ voffl = 1.944533E-8 minv = 0 nfactor = 0.583871
+ wnfactor = 4.630574E-8 eta0 = 9 etab = -2.1692E-4
+ dsub = 0.42 cit = 9.258412E-8 cdsc = 0
+ cdscb = 1.415095E-7 cdscd = 1.5E-5 pclm = 0.12036
+ wpclm = -2.853728E-8 pdiblc1 = 8.636946E-7 wpdiblc1 = 1.9429E-13
+ pdiblc2 = 2.202222E-4 wpdiblc2 = -2.004022E-10 pdiblcb = 0
+ drout = 0.133416 wdrout = -2.00803E-8 pscbe1 = 2.413849E8
+ wpscbe1 = 33.447131 pscbe2 = 2.610489E-9 wpscbe2 = 1.218446E-14
+ pvag = 4.541944 delta = 7E-3 fprout = 0
+ pdits = 2.202222E-4 wpdits = -2.004022E-10 pditsl = 0
+ pditsd = 0 lambda = 0 vtl = 0
+ lc = 5E-9 xn = 3 alpha0 = 2.136231E-6
+ walpha0 = -2.807635E-13 alpha1 = 8.04907E-2 walpha1 = 4.232495E-7
+ beta0 = 25.77902 wbeta0 = -1.100208E-6 aigbacc = 1
+ bigbacc = 0 cigbacc = 0 nigbacc = 1
+ aigbinv = 0.35 bigbinv = 0.03 cigbinv = 6E-3
+ eigbinv = 1.1 nigbinv = 3 aigc = 0.43
+ bigc = 0.054 cigc = 0.075 aigsd = 0.43
+ bigsd = 0.054 cigsd = 0.075 dlcig = 0
+ nigc = 1 poxedge = 1 pigcd = 1
+ ntox = 1 toxref = 1.16E-8 agidl = 0
+ bgidl = 2.3E9 cgidl = 0.5 egidl = 0.8
+ noia = 2.5E41 noib = 0 noic = 0
+ em = 4.1E7 af = 1 ef = 1
+ kf = 0 lintnoi = 0 tnoia = 7.6E6
+ tnoib = 7.2E6 ntnoi = 1 rnoia = 0.8
+ rnoib = 0.38 xpart = 0 cgso = {2.678273E-10/sw_func_tox_hv_ratio}
+ cgdo = {2.678273E-10/sw_func_tox_hv_ratio} cgbo = {0/sw_func_tox_hv_ratio} ckappas = 0.6
+ cf = 0 clc = 1E-7 cle = 0.6
+ dlc = 6.0712E-8 dwc = 0 vfbcv = -1
+ noff = 4 voffcv = 0.216 acde = 1.16
+ moin = 15 cgsl = {3.85585E-11/sw_func_tox_hv_ratio} cgdl = {3.85585E-11/sw_func_tox_hv_ratio}
+ ijthsrev = 0.1 ijthsfwd = 0.1 xjbvs = 1
+ bvs = 12.69 jss = 4.2966E-4 jsws = 8.04E-10
+ cjs = {8.310E-04*sw_func_nsd_pw_cj} mjs = 0.28329 mjsws = 0.057926
+ cjsws = {8.887314E-11*sw_func_nsd_pw_cj} cjswgs = {3.736446E-11*sw_func_nsd_pw_cj} mjswgs = 0.33
+ pbs = 0.66345 pbsws = 1 pbswgs = 0.2442
+ xrcrg1 = 12 xrcrg2 = 1 rbpb = 50
+ rbpd = 50 rbps = 50 rbdb = 50
+ rbsb = 50 gbmin = 1E-12 tnom = 30
+ ute = -1.464 kt1 = -0.37396 wkt1 = 7.334721E-9
+ kt1l = 0 kt2 = -0.01144 ua1 = 1E-9
+ ub1 = -7.128E-19 uc1 = 1E-11 at = 1.944108E4
+ wat = 4.649332E-4 prt = 0 njs = 1.5764
+ xtis = 0 tpb = 1.9685E-3 tpbsw = 1E-3
+ tpbswg = 0 tcj = 8.3E-4 tcjsw = 0
+ tcjswg = 0 tvoff = 0 tvfbsdoff = 0
+ saref = 2.54E-6 sbref = 2.54E-6 wlod = 0
+ ku0 = -3E-8 kvsat = 0.4 kvth0 = -7E-9
+ tku0 = 0 llodku0 = 0 wlodku0 = 1
+ llodvth = 0 wlodvth = 1 lku0 = 0
+ wku0 = 2E-7 pku0 = 0 lkvth0 = 0
+ wkvth0 = 8E-7 pkvth0 = 0 stk2 = 0
+ lodk2 = 1 steta0 = 0 lodeta0 = 1

.model nhvnative_model.11 nmos
+ level = 54 lmin = 8E-6 lmax = 2.525E-5 wmin = 4.2E-7
+ wmax = 1E-6 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 1.16E-8
+ toxm = 1.16E-8 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 1E23 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {4.5E-8+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {6.93E-8-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = -4.6E-9 dwb = 1.92E-9 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = 0.038459 lvth0 = 2.72244E-8
+ k1 = 0.364 k2 = 0.041446 lk2 = -1.271545E-8
+ k3 = 1.4 k3b = -0.58 w0 = 0
+ lpe0 = -1.236227E-14 lpeb = 0 vbm = -3
+ dvtp0 = 0 dvtp1 = 0 dvt0 = 5.7
+ dvt1 = 0.21851 dvt2 = 0.04 dvt0w = 7.7
+ dvt1w = 1.272E6 dvt2w = -0.032 vfbsdoff = 0
+ u0 = 4.45181E-2 lu0 = -2.145301E-9 ua = 1.096856E-9
+ lua = -2.413176E-17 ub = -1.500717E-19 lub = -1.033446E-24
+ uc = 1.9159E-11 ud = 0 up = 0
+ lp = 1 eu = 1.67 vsat = 7.5917E4
+ a0 = 1.387857 la0 = -1.035676E-5 ags = 2.90552E-2
+ lags = 3.780528E-6 b0 = 5.734E-8 b1 = 4.9905E-8
+ keta = -7.522213E-3 lketa = -1.067247E-7 a1 = 0
+ a2 = 0.962934 rdsw = 430 rdswmin = 0
+ rdw = 0 rdwmin = 0 rsw = 0
+ rswmin = 0 prwb = 0 prwg = 1E-12
+ wr = 1 voff = 0 voffl = 1.944533E-8
+ minv = 0 nfactor = 0.701166 lnfactor = -9.975764E-8
+ eta0 = 9 etab = -2.1692E-4 dsub = 0.42
+ cit = 9.258412E-8 cdsc = 0 cdscb = 1.415095E-7
+ cdscd = 1.5E-5 pclm = 0.089 pdiblc1 = 1.0772E-6
+ pdiblc2 = 5.1E-4 pdiblcb = 0 drout = 0.11135
+ pscbe1 = 2.7814E8 pscbe2 = 1.6E-8 pvag = 4.541944
+ delta = 7E-3 fprout = 0 pdits = -2.630332E-3
+ lpdits = 6.539373E-8 pditsl = 0 pditsd = 0
+ lambda = 0 vtl = 0 lc = 5E-9
+ xn = 3 alpha0 = 2.97923E-6 lalpha0 = -2.08346E-11
+ alpha1 = 0.5456 beta0 = 20.117451 lbeta0 = -8.73756E-6
+ aigbacc = 1 bigbacc = 0 cigbacc = 0
+ nigbacc = 1 aigbinv = 0.35 bigbinv = 0.03
+ cigbinv = 6E-3 eigbinv = 1.1 nigbinv = 3
+ aigc = 0.43 bigc = 0.054 cigc = 0.075
+ aigsd = 0.43 bigsd = 0.054 cigsd = 0.075
+ dlcig = 0 nigc = 1 poxedge = 1
+ pigcd = 1 ntox = 1 toxref = 1.16E-8
+ agidl = 0 bgidl = 2.3E9 cgidl = 0.5
+ egidl = 0.8 noia = 2.5E41 noib = 0
+ noic = 0 em = 4.1E7 af = 1
+ ef = 1 kf = 0 lintnoi = 0
+ tnoia = 7.6E6 tnoib = 7.2E6 ntnoi = 1
+ rnoia = 0.8 rnoib = 0.38 xpart = 0
+ cgso = {2.678273E-10/sw_func_tox_hv_ratio} cgdo = {2.678273E-10/sw_func_tox_hv_ratio} cgbo = {0/sw_func_tox_hv_ratio}
+ ckappas = 0.6 cf = 0 clc = 1E-7
+ cle = 0.6 dlc = 6.0712E-8 dwc = 0
+ vfbcv = -1 noff = 4 voffcv = 0.216
+ acde = 1.16 moin = 15 cgsl = {3.85585E-11/sw_func_tox_hv_ratio}
+ cgdl = {3.85585E-11/sw_func_tox_hv_ratio} ijthsrev = 0.1 ijthsfwd = 0.1
+ xjbvs = 1 bvs = 12.69 jss = 4.2966E-4
+ jsws = 8.04E-10 cjs = {8.310E-04*sw_func_nsd_pw_cj} mjs = 0.28329
+ mjsws = 0.057926 cjsws = {8.887314E-11*sw_func_nsd_pw_cj} cjswgs = {3.736446E-11*sw_func_nsd_pw_cj}
+ mjswgs = 0.33 pbs = 0.66345 pbsws = 1
+ pbswgs = 0.2442 xrcrg1 = 12 xrcrg2 = 1
+ rbpb = 50 rbpd = 50 rbps = 50
+ rbdb = 50 rbsb = 50 gbmin = 1E-12
+ tnom = 30 ute = -1.464 kt1 = -0.370524
+ lkt1 = 1.149679E-7 kt1l = 0 kt2 = -0.01144
+ ua1 = 1E-9 ub1 = -1.088076E-18 lub1 = 2.950191E-24
+ uc1 = 1E-11 at = 8.63772E4 lat = -0.496661
+ prt = 0 njs = 1.5764 xtis = 0
+ tpb = 1.9685E-3 tpbsw = 1E-3 tpbswg = 0
+ tcj = 8.3E-4 tcjsw = 0 tcjswg = 0
+ tvoff = 0 tvfbsdoff = 0 saref = 3E-6
+ sbref = 3E-6 wlod = 0 ku0 = -3E-8
+ kvsat = 0.4 kvth0 = -7E-9 tku0 = 0
+ llodku0 = 0 wlodku0 = 1 llodvth = 0
+ wlodvth = 1 lku0 = 0 wku0 = 2E-7
+ pku0 = 0 lkvth0 = 0 wkvth0 = 8E-7
+ pkvth0 = 0 stk2 = 0 lodk2 = 1
+ steta0 = 0 lodeta0 = 1

.model nhvnative_model.12 nmos
+ level = 54 lmin = 4E-6 lmax = 8E-6 wmin = 4.2E-7
+ wmax = 1E-6 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 1.16E-8
+ toxm = 1.16E-8 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 1E23 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {4.5E-8+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {6.93E-8-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = -4.6E-9 dwb = 1.92E-9 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = 4.57597E-2 lvth0 = -3.017008E-8
+ k1 = 0.364 k2 = 4.06964E-2 lk2 = -6.822741E-9
+ k3 = 1.4 k3b = -0.58 w0 = 0
+ lpe0 = -1.236227E-14 lpeb = 0 vbm = -3
+ dvtp0 = 0 dvtp1 = 0 dvt0 = 5.7
+ dvt1 = 0.21851 dvt2 = 0.04 dvt0w = 7.7
+ dvt1w = 1.272E6 dvt2w = -0.032 vfbsdoff = 0
+ u0 = 4.42452E-2 ua = 1.096187E-9 lua = -1.887385E-17
+ ub = -2.4364E-19 lub = -2.978683E-25 uc = 2.821794E-11
+ luc = -7.121596E-17 ud = 0 up = 0
+ lp = 1 eu = 1.67 vsat = 7.735441E4
+ lvsat = -0.0113 a0 = 4.41959E-2 la0 = 2.062916E-7
+ ags = 0.504411 lags = 4.356763E-8 b0 = 2.016994E-7
+ lb0 = -1.134867E-12 b1 = 4.9905E-8 keta = -0.021098
+ a1 = 0 a2 = 0.962934 rdsw = 430
+ rdswmin = 0 rdw = 0 rdwmin = 0
+ rsw = 0 rswmin = 0 prwb = 0
+ prwg = 1E-12 wr = 1 voff = 0
+ voffl = 1.944533E-8 minv = 0 nfactor = 0.690663
+ lnfactor = -1.718909E-8 eta0 = 9 etab = -2.1692E-4
+ dsub = 0.42 cit = 9.258412E-8 cdsc = 0
+ cdscb = 1.415095E-7 cdscd = 1.5E-5 pclm = 0.089
+ pdiblc1 = 1.0772E-6 pdiblc2 = 5.1E-4 pdiblcb = 0
+ drout = 0.11135 pscbe1 = 2.7814E8 pscbe2 = 1.6E-8
+ pvag = 4.541944 delta = 7E-3 fprout = 0
+ pdits = 5.688E-3 pditsl = 0 pditsd = 0
+ lambda = 0 vtl = 0 lc = 5E-9
+ xn = 3 alpha0 = 3.2899E-7 alpha1 = 0.5456
+ beta0 = 19.006 aigbacc = 1 bigbacc = 0
+ cigbacc = 0 nigbacc = 1 aigbinv = 0.35
+ bigbinv = 0.03 cigbinv = 6E-3 eigbinv = 1.1
+ nigbinv = 3 aigc = 0.43 bigc = 0.054
+ cigc = 0.075 aigsd = 0.43 bigsd = 0.054
+ cigsd = 0.075 dlcig = 0 nigc = 1
+ poxedge = 1 pigcd = 1 ntox = 1
+ toxref = 1.16E-8 agidl = 0 bgidl = 2.3E9
+ cgidl = 0.5 egidl = 0.8 noia = 2.5E41
+ noib = 0 noic = 0 em = 4.1E7
+ af = 1 ef = 1 kf = 0
+ lintnoi = 0 tnoia = 7.6E6 tnoib = 7.2E6
+ ntnoi = 1 rnoia = 0.8 rnoib = 0.38
+ xpart = 0 cgso = {2.678273E-10/sw_func_tox_hv_ratio} cgdo = {2.678273E-10/sw_func_tox_hv_ratio}
+ cgbo = {0/sw_func_tox_hv_ratio} ckappas = 0.6 cf = 0
+ clc = 1E-7 cle = 0.6 dlc = 6.0712E-8
+ dwc = 0 vfbcv = -1 noff = 4
+ voffcv = 0.216 acde = 1.16 moin = 15
+ cgsl = {3.85585E-11/sw_func_tox_hv_ratio} cgdl = {3.85585E-11/sw_func_tox_hv_ratio} ijthsrev = 0.1
+ ijthsfwd = 0.1 xjbvs = 1 bvs = 12.69
+ jss = 4.2966E-4 jsws = 8.04E-10 cjs = {8.310E-04*sw_func_nsd_pw_cj}
+ mjs = 0.28329 mjsws = 0.057926 cjsws = {8.887314E-11*sw_func_nsd_pw_cj}
+ cjswgs = {3.736446E-11*sw_func_nsd_pw_cj} mjswgs = 0.33 pbs = 0.66345
+ pbsws = 1 pbswgs = 0.2442 xrcrg1 = 12
+ xrcrg2 = 1 rbpb = 50 rbpd = 50
+ rbps = 50 rbdb = 50 rbsb = 50
+ gbmin = 1E-12 tnom = 30 ute = -1.464
+ kt1 = -0.356914 lkt1 = 7.968453E-9 kt1l = 0
+ kt2 = -0.01144 ua1 = 1E-9 ub1 = -7.128E-19
+ uc1 = 1E-11 at = 2.32E4 prt = 0
+ njs = 1.5764 xtis = 0 tpb = 1.9685E-3
+ tpbsw = 1E-3 tpbswg = 0 tcj = 8.3E-4
+ tcjsw = 0 tcjswg = 0 tvoff = 0
+ tvfbsdoff = 0 saref = 3E-6 sbref = 3E-6
+ wlod = 0 ku0 = -3E-8 kvsat = 0.4
+ kvth0 = -7E-9 tku0 = 0 llodku0 = 0
+ wlodku0 = 1 llodvth = 0 wlodvth = 1
+ lku0 = 0 wku0 = 2E-7 pku0 = 0
+ lkvth0 = 0 wkvth0 = 8E-7 pkvth0 = 0
+ stk2 = 0 lodk2 = 1 steta0 = 0
+ lodeta0 = 1

.model nhvnative_model.13 nmos
+ level = 54 lmin = 2E-6 lmax = 4E-6 wmin = 4.2E-7
+ wmax = 1E-6 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 1.16E-8
+ toxm = 1.16E-8 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 1E23 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {4.5E-8+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {6.93E-8-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = -4.6E-9 dwb = 1.92E-9 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = 4.69399E-2 lvth0 = -3.47273E-8
+ k1 = 0.364 k2 = 4.03756E-2 lk2 = -5.583946E-9
+ k3 = 1.4 k3b = -0.58 w0 = 0
+ lpe0 = -1.236227E-14 lpeb = 0 vbm = -3
+ dvtp0 = 0 dvtp1 = 0 dvt0 = 5.7
+ dvt1 = 0.21851 dvt2 = 0.04 dvt0w = 7.7
+ dvt1w = 1.272E6 dvt2w = -0.032 vfbsdoff = 0
+ u0 = 4.41235E-2 lu0 = 3.345832E-10 ua = 1.093895E-9
+ lua = -1.002312E-17 ub = -2.094124E-19 lub = -4.300347E-25
+ uc = 9.7749E-12 ud = 0 up = 0
+ lp = 1 eu = 1.67 vsat = 6.840451E4
+ lvsat = 2.32591E-2 a0 = 0.15654 la0 = -2.27513E-7
+ ags = 0.52853 lags = -4.956684E-8 b0 = -9.2201E-8
+ b1 = 4.9905E-8 keta = -0.021098 a1 = 0
+ a2 = 0.962934 rdsw = 430 rdswmin = 0
+ rdw = 0 rdwmin = 0 rsw = 0
+ rswmin = 0 prwb = 0 prwg = 1E-12
+ wr = 1 voff = 0 voffl = 1.944533E-8
+ minv = 0 nfactor = 0.712911 lnfactor = -1.030991E-7
+ eta0 = 9 etab = -2.1692E-4 dsub = 0.42
+ cit = 9.258412E-8 cdsc = 0 cdscb = 1.415095E-7
+ cdscd = 1.5E-5 pclm = 0.089 pdiblc1 = 1.0772E-6
+ pdiblc2 = 5.1E-4 pdiblcb = 0 drout = 0.11135
+ pscbe1 = 2.7814E8 pscbe2 = 1.6E-8 pvag = 4.541944
+ delta = 7E-3 fprout = 0 pdits = -3.723238E-3
+ lpdits = 3.634056E-8 pditsl = 0 pditsd = 0
+ lambda = 0 vtl = 0 lc = 5E-9
+ xn = 3 alpha0 = -1.065859E-6 lalpha0 = 5.386071E-12
+ alpha1 = 0.5456 beta0 = 16.126414 lbeta0 = 1.111923E-5
+ aigbacc = 1 bigbacc = 0 cigbacc = 0
+ nigbacc = 1 aigbinv = 0.35 bigbinv = 0.03
+ cigbinv = 6E-3 eigbinv = 1.1 nigbinv = 3
+ aigc = 0.43 bigc = 0.054 cigc = 0.075
+ aigsd = 0.43 bigsd = 0.054 cigsd = 0.075
+ dlcig = 0 nigc = 1 poxedge = 1
+ pigcd = 1 ntox = 1 toxref = 1.16E-8
+ agidl = 0 bgidl = 2.3E9 cgidl = 0.5
+ egidl = 0.8 noia = 2.5E41 noib = 0
+ noic = 0 em = 4.1E7 af = 1
+ ef = 1 kf = 0 lintnoi = 0
+ tnoia = 7.6E6 tnoib = 7.2E6 ntnoi = 1
+ rnoia = 0.8 rnoib = 0.38 xpart = 0
+ cgso = {2.678273E-10/sw_func_tox_hv_ratio} cgdo = {2.678273E-10/sw_func_tox_hv_ratio} cgbo = {0/sw_func_tox_hv_ratio}
+ ckappas = 0.6 cf = 0 clc = 1E-7
+ cle = 0.6 dlc = 6.0712E-8 dwc = 0
+ vfbcv = -1 noff = 4 voffcv = 0.216
+ acde = 1.16 moin = 15 cgsl = {3.85585E-11/sw_func_tox_hv_ratio}
+ cgdl = {3.85585E-11/sw_func_tox_hv_ratio} ijthsrev = 0.1 ijthsfwd = 0.1
+ xjbvs = 1 bvs = 12.69 jss = 4.2966E-4
+ jsws = 8.04E-10 cjs = {8.310E-04*sw_func_nsd_pw_cj} mjs = 0.28329
+ mjsws = 0.057926 cjsws = {8.887314E-11*sw_func_nsd_pw_cj} cjswgs = {3.736446E-11*sw_func_nsd_pw_cj}
+ mjswgs = 0.33 pbs = 0.66345 pbsws = 1
+ pbswgs = 0.2442 xrcrg1 = 12 xrcrg2 = 1
+ rbpb = 50 rbpd = 50 rbps = 50
+ rbdb = 50 rbsb = 50 gbmin = 1E-12
+ tnom = 30 ute = -1.464 kt1 = -0.344566
+ lkt1 = -3.971155E-8 kt1l = 0 kt2 = -0.01144
+ ua1 = 1E-9 ub1 = -7.128E-19 uc1 = 1E-11
+ at = 3.57235E4 lat = -4.83582E-2 prt = 0
+ njs = 1.5764 xtis = 0 tpb = 1.9685E-3
+ tpbsw = 1E-3 tpbswg = 0 tcj = 8.3E-4
+ tcjsw = 0 tcjswg = 0 tvoff = 0
+ tvfbsdoff = 0 saref = 3E-6 sbref = 3E-6
+ wlod = 0 ku0 = -3E-8 kvsat = 0.4
+ kvth0 = -7E-9 tku0 = 0 llodku0 = 0
+ wlodku0 = 1 llodvth = 0 wlodvth = 1
+ lku0 = 0 wku0 = 2E-7 pku0 = 0
+ lkvth0 = 0 wkvth0 = 8E-7 pkvth0 = 0
+ stk2 = 0 lodk2 = 1 steta0 = 0
+ lodeta0 = 1

.model nhvnative_model.14 nmos
+ level = 54 lmin = 1E-6 lmax = 2E-6 wmin = 4.2E-7
+ wmax = 1E-6 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 1.16E-8
+ toxm = 1.16E-8 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 1E23 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {4.5E-8+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {6.93E-8-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = -4.6E-9 dwb = 1.92E-9 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = -3.147271E-3 lvth0 = 5.850505E-8
+ wvth0 = 2.118442E-8 pvth0 = -3.943269E-14 k1 = 0.364
+ k2 = 0.038204 lk2 = -1.541833E-9 wk2 = -2.354143E-9
+ pk2 = 4.382002E-15 k3 = 1.4 k3b = -0.58
+ w0 = 0 lpe0 = -1.236227E-14 lpeb = 0
+ vbm = -3 dvtp0 = 0 dvtp1 = 0
+ dvt0 = 5.7 dvt1 = 0.21851 dvt2 = 0.04
+ dvt0w = 7.7 dvt1w = 1.272E6 dvt2w = -0.032
+ vfbsdoff = 0 u0 = 4.86391E-2 lu0 = -8.070886E-9
+ wu0 = -3.540505E-9 pu0 = 6.590296E-15 ua = 1.134458E-9
+ lua = -8.552674E-17 wua = -3.813589E-17 pua = 7.098614E-23
+ ub = -2.224612E-19 lub = -4.057457E-25 wub = -8.893186E-26
+ pub = 1.655378E-31 uc = 1.18829E-11 luc = -3.923829E-18
+ wuc = -1.918279E-18 puc = 3.570684E-24 ud = 0
+ up = 0 lp = 1 eu = 1.67
+ vsat = 8.688481E4 lvsat = -1.11401E-2 wvsat = -6.134024E-3
+ pvsat = 1.141787E-8 a0 = 3.572218E-3 la0 = 5.722089E-8
+ ags = 0.494607 lags = 1.357864E-8 b0 = -5.29454E-8
+ lb0 = -7.307038E-14 wb0 = -3.57226E-14 pb0 = 6.649404E-20
+ b1 = 5.071436E-8 lb1 = -1.506547E-15 wb1 = -7.365199E-16
+ pb1 = 1.370958E-21 keta = -2.98778E-2 lketa = 1.634267E-8
+ wketa = 7.989595E-9 pketa = -1.487183E-14 a1 = 0
+ a2 = 0.962934 rdsw = 430 rdswmin = 0
+ rdw = 0 rdwmin = 0 rsw = 0
+ rswmin = 0 prwb = 0 prwg = 1E-12
+ wr = 1 voff = 0 voffl = 1.944533E-8
+ minv = 0 nfactor = 0.684897 lnfactor = -5.095433E-8
+ wnfactor = -7.064686E-9 pnfactor = 1.315021E-14 eta0 = 9
+ etab = -2.1692E-4 dsub = 0.42 cit = 9.258412E-8
+ cdsc = 0 cdscb = 1.415095E-7 cdscd = 1.5E-5
+ pclm = 0.089 pdiblc1 = 1.0772E-6 pdiblc2 = 9.49314E-4
+ lpdiblc2 = -8.177391E-10 pdiblcb = 0 drout = 0.11135
+ pscbe1 = 2.7814E8 pscbe2 = 1.6E-8 pvag = 4.541944
+ delta = 7E-3 fprout = 0 pdits = 2.94101E-2
+ lpdits = -2.533388E-8 pditsl = 0 pditsd = 0
+ lambda = 0 vtl = 0 lc = 5E-9
+ xn = 3 alpha0 = 1.510454E-6 lalpha0 = 5.905221E-13
+ walpha0 = 2.88694E-13 palpha0 = -5.373751E-19 alpha1 = 0.417246
+ lalpha1 = 2.389183E-7 walpha1 = 1.168022E-7 palpha1 = -2.174157E-13
+ beta0 = 18.768149 lbeta0 = 6.201907E-6 wbeta0 = 1.095815E-6
+ pbeta0 = -2.039751E-12 aigbacc = 1 bigbacc = 0
+ cigbacc = 0 nigbacc = 1 aigbinv = 0.35
+ bigbinv = 0.03 cigbinv = 6E-3 eigbinv = 1.1
+ nigbinv = 3 aigc = 0.43 bigc = 0.054
+ cigc = 0.075 aigsd = 0.43 bigsd = 0.054
+ cigsd = 0.075 dlcig = 0 nigc = 1
+ poxedge = 1 pigcd = 1 ntox = 1
+ toxref = 1.16E-8 agidl = 0 bgidl = 2.3E9
+ cgidl = 0.5 egidl = 0.8 noia = 2.5E41
+ noib = 0 noic = 0 em = 4.1E7
+ af = 1 ef = 1 kf = 0
+ lintnoi = 0 tnoia = 7.6E6 tnoib = 7.2E6
+ ntnoi = 1 rnoia = 0.8 rnoib = 0.38
+ xpart = 0 cgso = {2.678273E-10/sw_func_tox_hv_ratio} cgdo = {2.678273E-10/sw_func_tox_hv_ratio}
+ cgbo = {0/sw_func_tox_hv_ratio} ckappas = 0.6 cf = 0
+ clc = 1E-7 cle = 0.6 dlc = 6.0712E-8
+ dwc = 0 vfbcv = -1 noff = 4
+ voffcv = 0.216 acde = 1.16 moin = 15
+ cgsl = {3.85585E-11/sw_func_tox_hv_ratio} cgdl = {3.85585E-11/sw_func_tox_hv_ratio} ijthsrev = 0.1
+ ijthsfwd = 0.1 xjbvs = 1 bvs = 12.69
+ jss = 4.2966E-4 jsws = 8.04E-10 cjs = {8.310E-04*sw_func_nsd_pw_cj}
+ mjs = 0.28329 mjsws = 0.057926 cjsws = {8.887314E-11*sw_func_nsd_pw_cj}
+ cjswgs = {3.736446E-11*sw_func_nsd_pw_cj} mjswgs = 0.33 pbs = 0.66345
+ pbsws = 1 pbswgs = 0.2442 xrcrg1 = 12
+ xrcrg2 = 1 rbpb = 50 rbpd = 50
+ rbps = 50 rbdb = 50 rbsb = 50
+ gbmin = 1E-12 tnom = 30 ute = -1.464
+ kt1 = -0.358725 lkt1 = -1.335585E-8 wkt1 = -6.5294E-9
+ pkt1 = 1.215383E-14 kt1l = 0 kt2 = -0.01144
+ ua1 = 1E-9 ub1 = -8.176045E-19 lub1 = 1.95083E-25
+ wub1 = 9.537206E-26 pub1 = -1.775255E-31 uc1 = 1E-11
+ at = 723.4192 lat = 1.67909E-2 wat = 2.069427E-4
+ pat = -3.852032E-10 prt = 0 njs = 1.5764
+ xtis = 0 tpb = 1.9685E-3 tpbsw = 1E-3
+ tpbswg = 0 tcj = 8.3E-4 tcjsw = 0
+ tcjswg = 0 tvoff = 0 tvfbsdoff = 0
+ saref = 3E-6 sbref = 3E-6 wlod = 0
+ ku0 = -3E-8 kvsat = 0.4 kvth0 = -7E-9
+ tku0 = 0 llodku0 = 0 wlodku0 = 1
+ llodvth = 0 wlodvth = 1 lku0 = 0
+ wku0 = 2E-7 pku0 = 0 lkvth0 = 0
+ wkvth0 = 8E-7 pkvth0 = 0 stk2 = 0
+ lodk2 = 1 steta0 = 0 lodeta0 = 1

.model nhvnative_model.15 nmos
+ level = 54 lmin = 9E-7 lmax = 1E-6 wmin = 4.2E-7
+ wmax = 1E-6 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 1.16E-8
+ toxm = 1.16E-8 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 1E23 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {4.5E-8+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {6.93E-8-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = -4.6E-9 dwb = 1.92E-9 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = 0.122908 lvth0 = -5.007906E-8
+ wvth0 = -7.749753E-8 pvth0 = 4.557195E-14 k1 = 0.364
+ k2 = 5.84719E-2 lk2 = -1.900056E-8 wk2 = -1.733964E-8
+ pk2 = 1.729051E-14 k3 = 1.4 k3b = -0.58
+ w0 = 0 lpe0 = -1.236227E-14 lpeb = 0
+ vbm = -3 dvtp0 = 0 dvtp1 = 0
+ dvt0 = 5.7 dvt1 = 0.21851 dvt2 = 0.04
+ dvt0w = 7.7 dvt1w = 1.272E6 dvt2w = -0.032
+ vfbsdoff = 0 u0 = 3.78825E-2 lu0 = 1.194882E-9
+ wu0 = 5.372472E-9 pu0 = -1.087343E-15 ua = 2.140063E-10
+ lua = 7.0735E-16 wua = 7.915305E-16 pua = -6.436885E-22
+ ub = 6.793519E-19 lub = -1.182567E-24 wub = -1.146047E-24
+ pub = 1.076136E-30 uc = -1.130509E-11 luc = 1.60503E-17
+ wuc = 1.918279E-17 puc = -1.460578E-23 ud = 0
+ up = 0 lp = 1 eu = 1.67
+ vsat = 4.773131E4 lvsat = 2.25867E-2 wvsat = 0.030982
+ pvsat = -2.05539E-8 a0 = 0.07 ags = 0.51037
+ b0 = -4.84757E-7 lb0 = 2.988922E-13 wb0 = 3.57226E-13
+ pb0 = -2.719919E-19 b1 = 4.181137E-8 lb1 = 6.162486E-15
+ wb1 = 7.365199E-15 pb1 = -5.607863E-21 keta = 7.18723E-2
+ lketa = -7.130483E-8 wketa = -8.460296E-8 pketa = 6.488739E-14
+ a1 = 0 a2 = 0.962934 rdsw = 430
+ rdswmin = 0 rdw = 0 rdwmin = 0
+ rsw = 0 rswmin = 0 prwb = 0
+ prwg = 1E-12 wr = 1 voff = 0
+ voffl = 1.944533E-8 minv = 0 nfactor = 0.499775
+ lnfactor = 1.085096E-7 wnfactor = 1.228331E-7 pnfactor = -9.874375E-14
+ eta0 = 9 etab = -2.1692E-4 dsub = 0.42
+ cit = 9.258412E-8 cdsc = 0 cdscb = 1.415095E-7
+ cdscd = 1.5E-5 pclm = 0.089 pdiblc1 = 1.0772E-6
+ pdiblc2 = 0 pdiblcb = 0 drout = 0.11135
+ pscbe1 = 2.7814E8 pscbe2 = 1.6E-8 pvag = 4.541944
+ delta = 7E-3 fprout = 0 pdits = 0
+ pditsl = 0 pditsd = 0 lambda = 0
+ vtl = 0 lc = 5E-9 xn = 3
+ alpha0 = 5.330268E-6 lalpha0 = -2.699866E-12 walpha0 = -3.187337E-12
+ palpha0 = 2.456878E-18 alpha1 = 1.829141 lalpha1 = -9.772881E-7
+ walpha1 = -1.168022E-6 palpha1 = 8.893322E-13 beta0 = 36.611926
+ lbeta0 = -9.168723E-6 wbeta0 = -1.095815E-5 pbeta0 = 8.343538E-12
+ aigbacc = 1 bigbacc = 0 cigbacc = 0
+ nigbacc = 1 aigbinv = 0.35 bigbinv = 0.03
+ cigbinv = 6E-3 eigbinv = 1.1 nigbinv = 3
+ aigc = 0.43 bigc = 0.054 cigc = 0.075
+ aigsd = 0.43 bigsd = 0.054 cigsd = 0.075
+ dlcig = 0 nigc = 1 poxedge = 1
+ pigcd = 1 ntox = 1 toxref = 1.16E-8
+ agidl = 0 bgidl = 2.3E9 cgidl = 0.5
+ egidl = 0.8 noia = 2.5E41 noib = 0
+ noic = 0 em = 4.1E7 af = 1
+ ef = 1 kf = 0 lintnoi = 0
+ tnoia = 7.6E6 tnoib = 7.2E6 ntnoi = 1
+ rnoia = 0.8 rnoib = 0.38 xpart = 0
+ cgso = {2.678273E-10/sw_func_tox_hv_ratio} cgdo = {2.678273E-10/sw_func_tox_hv_ratio} cgbo = {0/sw_func_tox_hv_ratio}
+ ckappas = 0.6 cf = 0 clc = 1E-7
+ cle = 0.6 dlc = 6.0712E-8 dwc = 0
+ vfbcv = -1 noff = 4 voffcv = 0.216
+ acde = 1.16 moin = 15 cgsl = {3.85585E-11/sw_func_tox_hv_ratio}
+ cgdl = {3.85585E-11/sw_func_tox_hv_ratio} ijthsrev = 0.1 ijthsfwd = 0.1
+ xjbvs = 1 bvs = 12.69 jss = 4.2966E-4
+ jsws = 8.04E-10 cjs = {8.310E-04*sw_func_nsd_pw_cj} mjs = 0.28329
+ mjsws = 0.057926 cjsws = {8.887314E-11*sw_func_nsd_pw_cj} cjswgs = {3.736446E-11*sw_func_nsd_pw_cj}
+ mjswgs = 0.33 pbs = 0.66345 pbsws = 1
+ pbswgs = 0.2442 xrcrg1 = 12 xrcrg2 = 1
+ rbpb = 50 rbpd = 50 rbps = 50
+ rbdb = 50 rbsb = 50 gbmin = 1E-12
+ tnom = 30 ute = -1.464 kt1 = -0.437652
+ lkt1 = 5.463171E-8 wkt1 = 6.5294E-8 pkt1 = -4.971485E-14
+ kt1l = 0 kt2 = -0.01144 ua1 = 1E-9
+ ub1 = 3.352446E-19 lub1 = -7.979811E-25 wub1 = -9.537206E-25
+ pub1 = 7.261628E-31 uc1 = 1E-11 at = 3.629677E4
+ lat = -0.013852 wat = -1.48737E-2 pat = 1.26053E-8
+ prt = 0 njs = 1.5764 xtis = 0
+ tpb = 1.9685E-3 tpbsw = 1E-3 tpbswg = 0
+ tcj = 8.3E-4 tcjsw = 0 tcjswg = 0
+ tvoff = 0 tvfbsdoff = 0 saref = 2.745E-6
+ sbref = 2.74E-6 wlod = 0 ku0 = -3E-8
+ kvsat = 0.4 kvth0 = -7E-9 tku0 = 0
+ llodku0 = 0 wlodku0 = 1 llodvth = 0
+ wlodvth = 1 lku0 = 0 wku0 = 2E-7
+ pku0 = 0 lkvth0 = 0 wkvth0 = 8E-7
+ pkvth0 = 0 stk2 = 0 lodk2 = 1
+ steta0 = 0 lodeta0 = 1
.ends sky130_fd_pr__nfet_05v0_nvt
