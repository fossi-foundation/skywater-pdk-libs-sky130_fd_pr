* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

******************************************************************
******************************************************************
*  *****************************************************
*  04/26/2021 Usman Suriono
*      Why     : New infrastructure of the sky130_fd_pr__pfet_01v8 20V model
*      What    : Converted from p20vhv1 models
*                Changed the parasitic Drain/Body diode from Deep Nwell-Sub to Pwell to
*                	Deep Nwell according to the device layout construction.
*                The device similar and correlated to sky130_fd_pr__pfet_g5v0d16v0.
*                Add "nf" (number of fingers)
*                Add process Monte Carlo
*                Changed the parasitic diode from internal dimension calculation
*                to receive it from PDK
*
*  *****************************************************
*
*  Pmos 20V VHV DE Model
*  -----------------------------------------------------

.subckt  sky130_fd_pr__pfet_20v0 d g s b  w=50u l=2u  nf=2   sa=0 sb=0 sd=0  mult=1
*** only estimated, the real values supplied and overwritten by PDK netlist
+ ad  = '9.73 * (w+11.72) - 5.75 * (w+6)'
+ pd  = '2 * ( 9.73 + 2*w + 11.72 + 5.75 + 6 )'
+ as  = '0.29  * w'
+ ps  = '2*(0.29 + w)'
*** preserve values, the resistance is dominated by "rldd" resistor
*** these values will be overwritten by PDK netlist
+ nrd = '0.205*nf/w'
+ nrs = '0.145*nf/w'


.param
+ sky130_fd_pr__pfet_20v0_agidl_diff  = 0
+ sky130_fd_pr__pfet_20v0_u0_diff     = -1.2404e-03
+ sky130_fd_pr__pfet_20v0_rdrift_mult = '9.1777e-01*1.05 * (sw_sky130_fd_pr__pfet_01v8_de_rd_mult*sw_pw_rs_mc**3)**0.7'


.param rdrift_tnom_sky130_fd_pr__pfet_20v0=1.595800e+004 vgdep=1.102900e-001 vth=7.000000e-001 vbdep=-5.260300e-001 
***** Swap these two lines if want to simulate in proplus
+ vth2=+1.048000e-001 hvvsat=1.878600e+000 avsat=7.467500e-001 
+ l_sky130_fd_pr__pfet_20v0=0.50 hvvbdep=-2.490600e-002 


.param tc1_rdrift_sky130_fd_pr__pfet_20v0=0.00621917042930238
.param tc2_rdrift_sky130_fd_pr__pfet_20v0=0.000021055807983754

.param
+rdrift_sky130_fd_pr__pfet_20v0='rdrift_tnom_sky130_fd_pr__pfet_20v0*((w-9.000000e-007)/w)*(1+tc1_rdrift_sky130_fd_pr__pfet_20v0*(temper-30)+tc2_rdrift_sky130_fd_pr__pfet_20v0*(temper-30)*(temper-30))*sky130_fd_pr__pfet_20v0_rdrift_mult'

****Zero out the drain diode params and put into seperate model
m1 d1 g s b sky130_fd_pr__pfet_20v0_base  w=w l=l_sky130_fd_pr__pfet_20v0 ad=0 as=as pd=0  ps=ps nrd=nrd nrs='nrs*sw_rdp/sw_pw_rs' nf=nf sa=sa sb=sb sd=sd
* + deltox  = 'sw_tox_hv_corner - sw_tox_hv_nom + sw_tox_hv_mc + sw_mm_tox_hv * mismatch_factor*MC_MM_SWITCH*AGAUSS(0,1.0,1)/sqrt(l_sky130_fd_pr__pfet_20v0*w*mult)'
+ delvto = '-0.0 + 1.52*sw_vth0_sky130_fd_pr__pfet_g5v0d16v0 +  sw_mm_vth0_sky130_fd_pr__pfet_g5v0d16v0 * mismatch_factor*MC_MM_SWITCH*AGAUSS(0,1.0,1)/sqrt(l_sky130_fd_pr__pfet_20v0*w*mult) + sw_vth0_sky130_fd_pr__pfet_g5v0d16v0_mc * 1.66'
* + mulu0   = sw_u0_sky130_fd_pr__pfet_g5v0d16v0
* + mulvsat = 'sw_vsat_sky130_fd_pr__pfet_g5v0d16v0**1.6'
* + delk1   = '-0.48*(sw_vth0_sky130_fd_pr__pfet_g5v0d16v0 + sw_vth0_sky130_fd_pr__pfet_g5v0d16v0_mc)'


rldd d d1 r='abs( (1/w)*(rdrift_sky130_fd_pr__pfet_20v0 /(1+0*(0-0-0 ))  )*  (1+0*pwr((abs(v(s,d)+vth2-min(v(s,d1),60))/(hvvsat*(1+hvvbdep*v(s,b)))),avsat)) )' tc1 = 0 tc2 = 0

xdnw1 d b sky130_fd_pr__model__parasitic__diode_pw2dn_defet area = {ad} perim = {pd} m = 0.5
xdnw2 d1 b sky130_fd_pr__model__parasitic__diode_pw2dn_defet area = {ad} perim = {pd} m = 0.5

****

.model sky130_fd_pr__pfet_20v0_base.0 pmos 
*
*DC IV MOS PARAMETERS
*
+ minr = 1e-6
+ lmin = 4.95e-07 lmax = 5.05e-07 wmin = 2.9995e-05 wmax = 1.0105e-03
+ level = 54
+ tnom = 30
+ version = 4.62
+ toxm = 1.175e-008
+ xj = 1.5e-007
+ lln = 1
+ lwn = 1
+ wln = 1
+ wwn = 1
+ lint = '4.5375e-08-sw_polycd'
+ ll = 0
+ lw = 0
+ lwl = 0
+ wint = '1.2277e-08+sw_activecd'
+ wl = 0
+ ww = 0
+ wwl = 0
+ xl = 0
+ xw = 0
+ mobmod = 0
+ binunit = 2
+ dwg = -4.7338e-009
+ dwb = 0
*NEW BSIM4 Parameters(Model Selectors)
+ igcmod = 0
+ igbmod = 0
+ rgatemod = 0
+ rbodymod = 1
+ trnqsmod = 0
+ acnqsmod = 0
+ fnoimod = 1
+ tnoimod = 1
+ permod = 1
+ geomod = 0
+ rdsmod = 0
+ tempmod = 0
*******
*NEW BSIM4 Parameters(4.4 Version)
+ lintnoi = 0
+ vfbsdoff = 0
+ lambda = 0
+ vtl = 0
+ lc = 5e-009
+ xn = 3
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
*NEW BSIM4 Parameters(Process Parameters)
+ epsrox = 3.9
+ toxe = 1.175e-08
+ dtox = 0
+ ndep = 1.7e+017
+ nsd = 1e+020
+ rshg = 0.1
****
+ rsh = {sw_pw_rs}
*
* THRESHOLD VOLTAGE PARAMETERS
*
+ vth0 = '-1.2314+8.3176e-02'
+ k1 = 0.66502
+ k2 = 0.038291
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300
+ dvt2w = 0
+ w0 = 0
+ k3b = -0.172
*NEW BSIM4 Parameters for Level 54
+ phin = 0
+ lpe0 = 0
+ lpeb = 0
+ vbm = -3
+ dvtp0 = 0
+ dvtp1 = 0
*
* MOBILITY PARAMETERS
*
+ vsat = 49870
+ ua = 2.1601000e-09
+ ub = 7.8839e-018
+ uc = -5.2815e-012
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.375
+ wr = 1
+ u0 = '0.020636+sky130_fd_pr__pfet_20v0_u0_diff'
+ a0 = 0.4683
+ keta = -0.15457
+ a1 = 0
+ a2 = 0.5
+ ags = 1.51
+ b0 = 0.0
+ b1 = 0.0
*NEW BSIM4 Parameters(Mobility Parameters)
+ eu = 1.67
+ rdswmin = 0
+ rdw = 0
+ rdwmin = 0
+ rsw = 0
+ rswmin = 0
*****
*
* SUBTHRESHOLD CURRENT PARAMETERS
*
+ voff = -0.10154
+ nfactor = 0.97411
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 5e-006
+ cdsc = 0
+ cdscb = 0
+ cdscd = 0
+ eta0 = 0.080055
+ etab = -0.0038503
+ dsub = 0.73391
*NEW BSIM4 Parameters(Sub-threshold parameters)
+ voffl = 0
+ minv = 0
*****
*
* ROUT PARAMETERS
*
+ pclm = 0.28871
+ pdiblc1 = 0.068215
+ pdiblc2 = 0
+ pdiblcb = -0.025
+ drout = 0.8996
+ pscbe1 = 6.0111000e+009
+ pscbe2 = 2.897300e-009
+ pvag = 0
+ delta = 0.01
+ alpha0 = 1.943700e-009
+ alpha1 = 0
+ beta0 = 87.25
*NEW BSIM4 Parameters(ROUT Parameters)
+ fprout = 0
+ pdits = 0
+ pditsl = 0
+ pditsd = 0
****
*NEW BSIM4 Parameters(GATE INDUCED DRAIN LEAKAGE MODEL PARAMTERS)
*****bgidl change on drain side, others copied from pfet
+ agidl = '1.3888e-08+sky130_fd_pr__pfet_20v0_agidl_diff'
+ bgidl = 1.16e+010
+ cgidl = 876
+ egidl = 0.66527
**************source side GIDL params copied from pfet
+ agisl = 1.3888e-08
+ bgisl = 1.6145e+009
+ cgisl = 876
+ egisl = 0.66527
****
****
*NEW BSIM4 Parameters(Gate Leakage Current Parameters)
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0
+ poxedge = 1
+ pigcd = 1
+ ntox = 1
+ toxref = 1.175e-008
*****
*
* TEMPERATURE EFFECTS PARAMETERS
*
+ kt1 = -0.61348
+ kt2 = -0.019032
+ at = 18000
+ ute = -1.3724
+ ua1 = 5.52e-010
+ ub1 = -2.16e-018
+ uc1 = -4.1496e-011
+ kt1l = 0
+ prt = 0
*NEW BSIM4 Parameters(HIGH SPEED RF MODEL PARAMETERS)
+ xrcrg1 = 12
+ xrcrg2 = 1
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ rbdb = 50
+ rbsb = 50
+ gbmin = 1e-012
****
*NEW BSIM4 Parameters(FLICKER and THERMAL NOISE PARAMETERS)
+ noia = 3.0000000E+40
+ noib = 8.5300000E+24
+ noic = 8.4000000E+07
+ em = 4.1000000E+07
+ af = 1
+ ef = 0.88
+ kf = 0
+ ntnoi = 1
*****
*NEW BSIM4 Parameters(LAYOUT DEPENDENT PARASITIC MODEL PARAMETERS)
+ dmcg = 0
+ dmcgt = 0
+ dmdg = 0
+ xgw = 0
+ xgl = 0
+ ngcon = 1
****
*
*DIODE DC IV PARAMTERS
*
*NEW BSIM4 Parameters(DIODE DC IV parameters)
+ diomod = 1
+ njs = 1.3632
+ jss = 2.1483e-05
+ jsws = 4.02e-12
+ xtis = 10
**+bvs        =        12.69
+ bvs = 24
+ xjbvs = 1
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
*
* DIODE and FET CAPACITANCE PARAMETERS
*
+ tpb = 0.001671
+ tpbsw = 0
+ tpbswg = 0
+ tcj = 0.00096
+ tcjsw = 3e-005
+ tcjswg = 0
+ cgdo = '3.50e-10 / sw_func_tox_hv_ratio'
+ cgso = '3.50e-10 / sw_func_tox_hv_ratio'
+ cgbo = 0
+ capmod = 2
+ xpart = 0
+ cgsl = '1.77e-11 / sw_func_tox_hv_ratio'
+ cgdl = '1.77e-11 / sw_func_tox_hv_ratio'
+ cf = 1.2e-011
+ clc = 1e-007
+ cle = 0.6
+ dlc = '-4.35e-07-sw_polycd'
+ dwc = {sw_activecd}
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4
+ voffcv = 0
+ ngate = 1e+023
+ lwc = 0
+ llc = 0
+ lwlc = 0
+ wlc = 0
+ wwc = 0
+ wwlc = 0
*NEW BSIM4 Parameters(FET and DIODE capacitance parameters)
+ ckappas = 0.6
+ cjs = '7.682E-04*sw_func_psd_nw_cj'
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = '9.9605453e-11*sw_func_psd_nw_cj'
+ mjsws = 0.24676
+ pbsws = 1
+ cjswgs = '1.47314e-10*sw_func_nsd_pw_cj'
+ mjswgs = 0.81
+ pbswgs = 3
*
*STRESS PARAMETERS
*
+ saref = 1.81e-06
+ sbref = 1.81e-06
+ wlod = 0.0
+ kvth0 = 3.5e-08
+ lkvth0 = 0.0
+ wkvth0 = 6.5e-07
+ pkvth0 = 0
+ llodvth = 0
+ wlodvth = 1
+ stk2 = 0
+ lodk2 = 1
+ lodeta0 = 1
+ ku0 = 7.0e-08
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0
+ llodku0 = 0
+ wlodku0 = 1
+ kvsat = 0.4
+ steta0 = 0
+ tku0 = 0
******

.ends sky130_fd_pr__pfet_20v0
*[Instances section]

*[analysis and output]

*simulator lang = spectre insensitive=yes

*simulator lang = spice
*[netlist end]

*.END
**** ; $&%*(C)Proplus Inc. All rights Reserved.
