* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

******************************************************************
******************************************************************
*  *****************************************************
*  04/24/2021 Usman Suriono
*      Why     : New scalable sky130_fd_pr__pfet_01v8 model
*      What    : Converted from discrete pshort model
*                Replaced rsh from 1 to calculated rsh from the original model.
*                PDK netlist nrd/nrs = ratio of distance the middle of the contact to Gate.
*
*  *****************************************************
*
*  Pmos Model
*  -----------------------------------------------------

.subckt  sky130_fd_pr__pfet_01v8  d g s b  mult=1
+ 
.param  l = 1 w = 1 nf = 1 ad = 0 as = 0 pd = 0 ps = 0 nrd = {0.14/w} nrs = {0.14/w} sa = 0 sb = 0 sd = 0
+ swx_nrds = {361*nf/w+1489}

Msky130_fd_pr__pfet_01v8  d g s b pshort_model l = {l} w = {w} ad = {ad} as = {as} pd = {pd} ps = {ps} nrd = {nrd} nrs = {nrs} sa = {sa} sb = {sb} sd = {sd} nf = {nf}
* + deltox = 0.3*(sw_tox_lv_corner - sw_tox_lv_nom) + sw_tox_lv_mc + sw_mm_tox_lv * mismatch_factor*MC_MM_SWITCH*AGAUSS(0,1.0,1)/sqrt(l*w*mult)
+ delvto = {(sw_vth0_sky130_fd_pr__pfet_01v8+sw_vth0_sky130_fd_pr__pfet_01v8_mc)*(0.0230*8/l+0.9770)*(0.028*7/w+0.972)*(0.0005*56/(w*l)+0.9995)+sw_mm_vth0_sky130_fd_pr__pfet_01v8*mismatch_factor*MC_MM_SWITCH*AGAUSS(0,1.0,1)/sqrt(l*w*mult)}
* + mulu0  = sw_u0_sky130_fd_pr__pfet_01v8
* + mulvsat= sw_vsat_sky130_fd_pr__pfet_01v8



.model pshort_model.1 pmos
+ level = 54 lmin = 8E-6 lmax = 2.02E-5 wmin = 7E-6
+ wmax = 1.01E-3 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 4.23E-9
+ toxm = 4.23E-9 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 9.999999999999999E22 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {7.3039E-9+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {-1.3994E-8-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = -5.722E-9 dwb = -1.7864E-8 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = -1.05955351 k1 = 0.43448553
+ k2 = 0.019777346 k3 = -15.845 k3b = 2
+ w0 = 0 lpe0 = 0 lpeb = 0
+ vbm = -3 dvtp0 = 0 dvtp1 = 0
+ dvt0 = 4.4955 dvt1 = 0.294 dvt2 = 0.015
+ dvt0w = -4.9772 dvt1w = 1.1472E6 dvt2w = -8.96E-3
+ vfbsdoff = 0 u0 = 0.0104766 ua = -5.6585471E-10
+ ub = 9.3302446E-19 uc = -6.6549964E-11 ud = 0
+ up = 0 lp = 1 eu = 1.67
+ vsat = 1.603125E5 a0 = 1.23682 ags = 0.2261248
+ b0 = 0 b1 = 0 keta = 5.1290095E-3
+ a1 = 0 a2 = 0.9995 rdsw = 547.88
+ rdswmin = 0 rdw = 0 rdwmin = 0
+ rsw = 0 rswmin = 0 prwb = -0.32348
+ prwg = 0.1376 wr = 1 voff = -0.25706245
+ voffl = 0 minv = 0 nfactor = 1.3376708
+ eta0 = 0.08 etab = -0.07 dsub = 0.56
+ cit = 1E-5 cdsc = 1.3E-4 cdscb = 7.8E-4
+ cdscd = 0 pclm = 1.5228006E-3 pdiblc1 = 0.39
+ pdiblc2 = 2.9632464E-3 pdiblcb = -0.025 drout = 0.56
+ pscbe1 = 8E8 pscbe2 = 9.3760948E-9 pvag = 0
+ delta = 0.01 fprout = 0 pdits = 0
+ pditsl = 0 pditsd = 0 lambda = 0
+ vtl = 0 lc = 5E-9 xn = 3
+ alpha0 = 1E-10 alpha1 = 1E-10 beta0 = 4.6464006
+ aigbacc = 0.43 bigbacc = 0.054 cigbacc = 0.075
+ nigbacc = 1 aigbinv = 0.35 bigbinv = 0.03
+ cigbinv = 6E-3 eigbinv = 1.1 nigbinv = 3
+ aigc = 0.43 bigc = 0.054 cigc = 0.075
+ aigsd = 0.43 bigsd = 0.054 cigsd = 0.075
+ dlcig = 0 nigc = 1 poxedge = 1
+ pigcd = 1 ntox = 1 toxref = 4.23E-9
+ agidl = 1E-10 bgidl = 1.181082E9 cgidl = 300
+ egidl = 0.1 noia = 1.5E42 noib = 0
+ noic = 0 em = 4.1E7 af = 1
+ ef = 1 kf = 0 lintnoi = -2E-7
+ tnoia = 2.5E7 tnoib = 0 ntnoi = 1
+ rnoia = 0.69 rnoib = 0.34 xpart = 0
+ cgso = {5.248925E-11/sw_func_tox_lv_ratio} cgdo = {5.248925E-11/sw_func_tox_lv_ratio} cgbo = {0/sw_func_tox_lv_ratio}
+ ckappas = 0.6 cf = 1.2E-11 clc = 1E-7
+ cle = 0.6 dlc = -3E-9 dwc = 0
+ vfbcv = -0.14469 noff = 3.9 voffcv = -0.10701
+ acde = 0.8 moin = 18.13 cgsl = {9.548271750000001E-12/sw_func_tox_lv_ratio}
+ cgdl = {9.548271750000001E-12/sw_func_tox_lv_ratio} ijthsrev = 0.1 ijthsfwd = 0.1
+ xjbvs = 1 bvs = 12.69 jss = 2.1483E-5
+ jsws = 8.040000000000001E-10 cjs = {sw_psd_nw_cj} mjs = 0.34629
+ mjsws = 0.29781 cjsws = {9.888891999999999E-11*sw_func_psd_nw_cj} cjswgs = {2.39155046E-10*sw_func_psd_nw_cj}
+ mjswgs = 0.9274 pbs = 0.6587 pbsws = 0.7418
+ pbswgs = 1.4338 xrcrg1 = 12 xrcrg2 = 1
+ rbpb = 50 rbpd = 50 rbps = 50
+ rbdb = 50 rbsb = 50 gbmin = 1E-12
+ tnom = 30 ute = -0.33954 kt1 = -0.4485
+ kt1l = 0 kt2 = -7.5706E-3 ua1 = 1.6104E-9
+ ub1 = -5.609E-19 uc1 = -1.0858E-10 at = 9.09E4
+ prt = 0 njs = 1.3632 xtis = 5.2
+ tpb = 2.0386E-3 tpbsw = 1.246E-3 tpbswg = 0
+ tcj = 1.2407E-3 tcjsw = 3.7357E-4 tcjswg = 2E-12
+ tvoff = 0 tvfbsdoff = 0 saref = 3E-6
+ sbref = 3E-6 wlod = 0 ku0 = 4.5E-8
+ kvsat = 0.5 kvth0 = 3.29E-8 tku0 = 0
+ llodku0 = 0 wlodku0 = 1 llodvth = 0
+ wlodvth = 1 lku0 = 0 wku0 = 2.5E-7
+ pku0 = 0 lkvth0 = 0 wkvth0 = 2E-7
+ pkvth0 = 0 stk2 = 0 lodk2 = 1
+ steta0 = 0 lodeta0 = 1

.model pshort_model.2 pmos
+ level = 54 lmin = 4E-6 lmax = 8E-6 wmin = 7E-6
+ wmax = 1.01E-3 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 4.23E-9
+ toxm = 4.23E-9 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 9.999999999999999E22 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {7.3039E-9+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {-1.3994E-8-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = -5.722E-9 dwb = -1.7864E-8 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = -1.06313713036384 lvth0 = 2.876926127746328E-8
+ k1 = 0.43813350754211 lk1 = -2.92859199323287E-8 k2 = 0.018505134186116
+ lk2 = 1.021330117531898E-8 k3 = -15.845 k3b = 2
+ w0 = 0 lpe0 = 0 lpeb = 0
+ vbm = -3 dvtp0 = 0 dvtp1 = 0
+ dvt0 = 4.4955 dvt1 = 0.294 dvt2 = 0.015
+ dvt0w = -4.9772 dvt1w = 1.1472E6 dvt2w = -8.96E-3
+ vfbsdoff = 0 u0 = 0.0102870831646 lu0 = 1.521438880389171E-9
+ ua = -5.773510610405899E-10 lua = 9.229256819764354E-17 ub = 9.280149419541299E-19
+ lub = 4.021635075802814E-26 uc = -7.3225399476844E-11 luc = 5.359031590287793E-17
+ ud = 0 up = 0 lp = 1
+ eu = 1.67 vsat = 2.67935304375E5 lvsat = -0.863994582048848
+ a0 = 1.328853483818 la0 = -7.38843703689098E-7 ags = 0.15379317220712
+ lags = 5.806774399417075E-7 b0 = 0 b1 = 0
+ keta = 0.021456825908407 lketa = -1.310795141928905E-7 a1 = 0
+ a2 = 1.2003959015 la2 = -1.612789886491182E-6 rdsw = 547.88
+ rdswmin = 0 rdw = 0 rdwmin = 0
+ rsw = 0 rswmin = 0 prwb = -0.32348
+ prwg = 0.1376 wr = 1 voff = -0.26700524634887
+ lvoff = 7.982064977517224E-8 voffl = 0 minv = 0
+ nfactor = 1.1833079277709 lnfactor = 1.239223285900749E-6 eta0 = 0.08
+ etab = -0.07 dsub = 0.56 cit = 1E-5
+ cdsc = 1.3E-4 cdscb = 7.8E-4 cdscd = 0
+ pclm = -0.433600672985592 lpclm = 3.493166024463448E-6 pdiblc1 = 0.39
+ pdiblc2 = 5.78918120501261E-3 lpdiblc2 = -2.268657070342358E-8 pdiblcb = -0.025
+ drout = 0.56 pscbe1 = 8E8 pscbe2 = 1.01417218694784E-8
+ lpscbe2 = -6.146444926247763E-15 pvag = 0 delta = 0.01
+ fprout = 0 pdits = 0 pditsl = 0
+ pditsd = 0 lambda = 0 vtl = 0
+ lc = 5E-9 xn = 3 alpha0 = 1E-10
+ alpha1 = 1E-10 beta0 = 3.2444736759574 lbeta0 = 1.12546525230909E-5
+ aigbacc = 0.43 bigbacc = 0.054 cigbacc = 0.075
+ nigbacc = 1 aigbinv = 0.35 bigbinv = 0.03
+ cigbinv = 6E-3 eigbinv = 1.1 nigbinv = 3
+ aigc = 0.43 bigc = 0.054 cigc = 0.075
+ aigsd = 0.43 bigsd = 0.054 cigsd = 0.075
+ dlcig = 0 nigc = 1 poxedge = 1
+ pigcd = 1 ntox = 1 toxref = 4.23E-9
+ agidl = 8.426709174077001E-11 lagidl = 1.263035987101993E-16 bgidl = 1.363431030754E9
+ lbgidl = -1.463895830704743E3 cgidl = 300 egidl = 0.1
+ noia = 1.5E42 noib = 0 noic = 0
+ em = 4.1E7 af = 1 ef = 1
+ kf = 0 lintnoi = -2E-7 tnoia = 2.5E7
+ tnoib = 0 ntnoi = 1 rnoia = 0.69
+ rnoib = 0.34 xpart = 0 cgso = {5.248925E-11/sw_func_tox_lv_ratio}
+ cgdo = {5.248925E-11/sw_func_tox_lv_ratio} cgbo = {0/sw_func_tox_lv_ratio} ckappas = 0.6
+ cf = 1.2E-11 clc = 1E-7 cle = 0.6
+ dlc = -3E-9 dwc = 0 vfbcv = -0.14469
+ noff = 3.9 voffcv = -0.10701 acde = 0.8
+ moin = 18.13 cgsl = {9.548271750000001E-12/sw_func_tox_lv_ratio} cgdl = {9.548271750000001E-12/sw_func_tox_lv_ratio}
+ ijthsrev = 0.1 ijthsfwd = 0.1 xjbvs = 1
+ bvs = 12.69 jss = 2.1483E-5 jsws = 8.040000000000001E-10
+ cjs = {sw_psd_nw_cj} mjs = 0.34629 mjsws = 0.29781
+ cjsws = {9.888891999999999E-11*sw_func_psd_nw_cj} cjswgs = {2.39155046E-10*sw_func_psd_nw_cj} mjswgs = 0.9274
+ pbs = 0.6587 pbsws = 0.7418 pbswgs = 1.4338
+ xrcrg1 = 12 xrcrg2 = 1 rbpb = 50
+ rbpd = 50 rbps = 50 rbdb = 50
+ rbsb = 50 gbmin = 1E-12 tnom = 30
+ ute = -0.47442366324068 lute = 1.08284442989222E-6 kt1 = -0.43157364924622
+ lkt1 = -1.358845407351367E-7 kt1l = 0 kt2 = 9.803815075927001E-3
+ lkt2 = -1.39481595736561E-7 ua1 = 1.2238699414329E-9 lua1 = 3.103058671815977E-15
+ ub1 = -2.993962520201601E-19 lub1 = -2.099348950737179E-24 uc1 = -8.830298756835999E-11
+ luc1 = -1.627836124770568E-16 at = 8.786010766631E4 lat = 0.024404219176155
+ prt = 0 njs = 1.3632 xtis = 5.2
+ tpb = 2.0386E-3 tpbsw = 1.246E-3 tpbswg = 0
+ tcj = 1.2407E-3 tcjsw = 3.7357E-4 tcjswg = 2E-12
+ tvoff = 0 tvfbsdoff = 0 saref = 3E-6
+ sbref = 3E-6 wlod = 0 ku0 = 4.5E-8
+ kvsat = 0.5 kvth0 = 3.29E-8 tku0 = 0
+ llodku0 = 0 wlodku0 = 1 llodvth = 0
+ wlodvth = 1 lku0 = 0 wku0 = 2.5E-7
+ pku0 = 0 lkvth0 = 0 wkvth0 = 2E-7
+ pkvth0 = 0 stk2 = 0 lodk2 = 1
+ steta0 = 0 lodeta0 = 1

.model pshort_model.3 pmos
+ level = 54 lmin = 2E-6 lmax = 4E-6 wmin = 7E-6
+ wmax = 1.01E-3 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 4.23E-9
+ toxm = 4.23E-9 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 9.999999999999999E22 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {7.3039E-9+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {-1.3994E-8-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = -5.722E-9 dwb = -1.7864E-8 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = -1.06465013124466 lvth0 = 3.486361066939505E-8
+ k1 = 0.4242721924985 lk1 = 2.654729072755209E-8 k2 = 0.023299152360404
+ lk2 = -9.096946502494982E-9 k3 = -15.845 k3b = 2
+ w0 = 0 lpe0 = 0 lpeb = 0
+ vbm = -3 dvtp0 = 0 dvtp1 = 0
+ dvt0 = 4.4955 dvt1 = 0.294 dvt2 = 0.015
+ dvt0w = -4.9772 dvt1w = 1.1472E6 dvt2w = -8.96E-3
+ vfbsdoff = 0 u0 = 0.0121663223152 lu0 = -6.048113867357822E-9
+ ua = -2.310026979311001E-10 lua = -1.302794482227024E-15 ub = 7.527581526871801E-19
+ lub = 7.461485948438308E-25 uc = -8.0891709259708E-11 luc = 8.447011971253669E-17
+ ud = 0 up = 0 lp = 1
+ eu = 1.67 vsat = 5.34375E4 a0 = 1.171646870846
+ la0 = -1.056173531172382E-7 ags = 0.09441453032174 lags = 8.198538969123151E-7
+ b0 = 0 b1 = 0 keta = -5.464761922144001E-3
+ lketa = -2.263968147048703E-8 a1 = 0 a2 = 0.8
+ rdsw = 547.88 rdswmin = 0 rdw = 0
+ rdwmin = 0 rsw = 0 rswmin = 0
+ prwb = -0.32348 prwg = 0.1376 wr = 1
+ voff = -0.25410325634546 lvoff = 2.785158886531673E-8 voffl = 0
+ minv = 0 nfactor = 1.514261668126 lnfactor = -9.385440880471083E-8
+ eta0 = 0.160612523 leta0 = -3.24706275293724E-7 etab = -0.140472582563983
+ letab = 2.838627168967311E-7 dsub = 0.8641982 ldsub = -1.2253066992216E-6
+ cit = 1E-5 cdsc = 1.3E-4 cdscb = 7.8E-4
+ cdscd = 0 pclm = 0.46461195637154 lpclm = -1.248236680355267E-7
+ pdiblc1 = 0.39 pdiblc2 = -2.158869170793999E-5 lpdiblc2 = 7.191407113280418E-10
+ pdiblcb = -0.025 drout = 0.56 pscbe1 = 8E8
+ pscbe2 = 8.286433932649798E-9 lpscbe2 = 1.326632619842603E-15 pvag = 0
+ delta = 0.01 fprout = 0 pdits = 0
+ pditsl = 0 pditsd = 0 lambda = 0
+ vtl = 0 lc = 5E-9 xn = 3
+ alpha0 = 1E-10 alpha1 = 1E-10 beta0 = 3.8949963916396
+ lbeta0 = 8.63435483059559E-6 aigbacc = 0.43 bigbacc = 0.054
+ cigbacc = 0.075 nigbacc = 1 aigbinv = 0.35
+ bigbinv = 0.03 cigbinv = 6E-3 eigbinv = 1.1
+ nigbinv = 3 aigc = 0.43 bigc = 0.054
+ cigc = 0.075 aigsd = 0.43 bigsd = 0.054
+ cigsd = 0.075 dlcig = 0 nigc = 1
+ poxedge = 1 pigcd = 1 ntox = 1
+ toxref = 4.23E-9 agidl = 1.3146581651846E-10 lagidl = -6.381229830963865E-17
+ bgidl = 9.172524112336E8 lbgidl = 333.306294579994 cgidl = 300
+ egidl = 0.1 noia = 1.5E42 noib = 0
+ noic = 0 em = 4.1E7 af = 1
+ ef = 1 kf = 0 lintnoi = -2E-7
+ tnoia = 2.5E7 tnoib = 0 ntnoi = 1
+ rnoia = 0.69 rnoib = 0.34 xpart = 0
+ cgso = {5.248925E-11/sw_func_tox_lv_ratio} cgdo = {5.248925E-11/sw_func_tox_lv_ratio} cgbo = {0/sw_func_tox_lv_ratio}
+ ckappas = 0.6 cf = 1.2E-11 clc = 1E-7
+ cle = 0.6 dlc = -3E-9 dwc = 0
+ vfbcv = -0.14469 noff = 3.9 voffcv = -0.10701
+ acde = 0.8 moin = 18.13 cgsl = {9.548271750000001E-12/sw_func_tox_lv_ratio}
+ cgdl = {9.548271750000001E-12/sw_func_tox_lv_ratio} ijthsrev = 0.1 ijthsfwd = 0.1
+ xjbvs = 1 bvs = 12.69 jss = 2.1483E-5
+ jsws = 8.040000000000001E-10 cjs = {sw_psd_nw_cj} mjs = 0.34629
+ mjsws = 0.29781 cjsws = {9.888891999999999E-11*sw_func_psd_nw_cj} cjswgs = {2.39155046E-10*sw_func_psd_nw_cj}
+ mjswgs = 0.9274 pbs = 0.6587 pbsws = 0.7418
+ pbswgs = 1.4338 xrcrg1 = 12 xrcrg2 = 1
+ rbpb = 50 rbpd = 50 rbps = 50
+ rbdb = 50 rbsb = 50 gbmin = 1E-12
+ tnom = 30 ute = -0.17571011240618 lute = -1.203701683065358E-7
+ kt1 = -0.46636744099546 lkt1 = 4.264434905300925E-9 kt1l = 0
+ kt2 = -5.478318739885996E-3 lkt2 = -7.792534411207208E-8 ua1 = 2.345249984031E-9
+ lua1 = -1.41384668320866E-15 ub1 = -1.03151249939108E-18 lub1 = 8.496065082779174E-25
+ uc1 = -2.42518521215026E-10 luc1 = 4.583947064653101E-16 at = 1.07038244165516E5
+ lat = -0.052845084505008 prt = 0 njs = 1.3632
+ xtis = 5.2 tpb = 2.0386E-3 tpbsw = 1.246E-3
+ tpbswg = 0 tcj = 1.2407E-3 tcjsw = 3.7357E-4
+ tcjswg = 2E-12 tvoff = 0 tvfbsdoff = 0
+ saref = 3E-6 sbref = 3E-6 wlod = 0
+ ku0 = 4.5E-8 kvsat = 0.5 kvth0 = 3.29E-8
+ tku0 = 0 llodku0 = 0 wlodku0 = 1
+ llodvth = 0 wlodvth = 1 lku0 = 0
+ wku0 = 2.5E-7 pku0 = 0 lkvth0 = 0
+ wkvth0 = 2E-7 pkvth0 = 0 stk2 = 0
+ lodk2 = 1 steta0 = 0 lodeta0 = 1

.model pshort_model.4 pmos
+ level = 54 lmin = 1E-6 lmax = 2E-6 wmin = 7E-6
+ wmax = 1.01E-3 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 4.23E-9
+ toxm = 4.23E-9 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 9.999999999999999E22 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {7.3039E-9+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {-1.3994E-8-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = -5.722E-9 dwb = -1.7864E-8 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = -1.0639711628476 lvth0 = 3.34866709077786E-8
+ k1 = 0.354542539783 lk1 = 1.679581896787533E-7 k2 = 0.051575195178736
+ lk2 = -6.644042202555847E-8 k3 = -15.845 k3b = 2
+ w0 = 0 lpe0 = 0 lpeb = 0
+ vbm = -3 dvtp0 = 0 dvtp1 = 0
+ dvt0 = 4.4955 dvt1 = 0.294 dvt2 = 0.015
+ dvt0w = -4.9772 dvt1w = 1.1472E6 dvt2w = -8.96E-3
+ vfbsdoff = 0 u0 = 9.785784175199999E-3 lu0 = -1.220411085895497E-9
+ ua = -7.482355275187199E-10 lua = -2.538525106172862E-16 ub = 1.05727653665008E-18
+ lub = 1.285889663876778E-25 uc = -4.298706539394E-11 luc = 7.599956808485589E-18
+ ud = 0 up = 0 lp = 1
+ eu = 1.67 vsat = 3.512646375E4 lvsat = 0.037134561782565
+ a0 = 1.293787322276 la0 = -3.533167229318607E-7 ags = 0.3713411399114
+ lags = 2.582500557837996E-7 b0 = 0 b1 = 0
+ keta = -6.680825932651995E-3 lketa = -2.017351824994494E-8 a1 = 0
+ a2 = 0.6972012 la2 = 2.084747328143999E-7 rdsw = 547.88
+ rdswmin = 0 rdw = 0 rdwmin = 0
+ rsw = 0 rswmin = 0 prwb = -0.32348
+ prwg = 0.1376 wr = 1 voff = -0.2479929006116
+ lvoff = 1.545986076131745E-8 voffl = 0 minv = 0
+ nfactor = 1.2665691307516 lnfactor = 4.084630846801242E-7 eta0 = -0.502700126
+ leta0 = 1.020483817126488E-6 etab = 7.645320704060766 letab = -1.550563263885882E-5
+ dsub = 0.26 cit = 1E-5 cdsc = 1.3E-4
+ cdscb = 7.8E-4 cdscd = 0 pclm = 0.18260436541916
+ lpclm = 4.470843423248086E-7 pdiblc1 = 0.40860196713388 lpdiblc1 = -3.772456612390311E-8
+ pdiblc2 = 2.3332426360864E-4 lpdiblc2 = 2.021802969014813E-10 pdiblcb = -0.049934208571322
+ lpdiblcb = 5.0566275772138E-8 drout = 0.40005836936472 ldrout = 3.243597076287802E-7
+ pscbe1 = 7.9955987E8 pscbe2 = 8.9405959E-9 pvag = 0
+ delta = 0.01 fprout = 0 pdits = 0
+ pditsl = 0 pditsd = 0 lambda = 0
+ vtl = 0 lc = 5E-9 xn = 3
+ alpha0 = -4.5896723869156E-5 lalpha0 = 9.307820804476194E-11 alpha1 = 2.027988E-10
+ lalpha1 = -2.084747328144E-16 beta0 = -14.198337403152 lbeta0 = 4.532741864642742E-5
+ aigbacc = 0.43 bigbacc = 0.054 cigbacc = 0.075
+ nigbacc = 1 aigbinv = 0.35 bigbinv = 0.03
+ cigbinv = 6E-3 eigbinv = 1.1 nigbinv = 3
+ aigc = 0.43 bigc = 0.054 cigc = 0.075
+ aigsd = 0.43 bigsd = 0.054 cigsd = 0.075
+ dlcig = 0 nigc = 1 poxedge = 1
+ pigcd = 1 ntox = 1 toxref = 4.23E-9
+ agidl = 1E-10 bgidl = 7.978149151704E8 lbgidl = 575.5241033462108
+ cgidl = 300 egidl = 0.1 noia = 1.5E42
+ noib = 0 noic = 0 em = 4.1E7
+ af = 1 ef = 1 kf = 0
+ lintnoi = -2E-7 tnoia = 2.5E7 tnoib = 0
+ ntnoi = 1 rnoia = 0.69 rnoib = 0.34
+ xpart = 0 cgso = {5.248925E-11/sw_func_tox_lv_ratio} cgdo = {5.248925E-11/sw_func_tox_lv_ratio}
+ cgbo = {0/sw_func_tox_lv_ratio} ckappas = 0.6 cf = 1.2E-11
+ clc = 1E-7 cle = 0.6 dlc = -3E-9
+ dwc = 0 vfbcv = -0.14469 noff = 3.9
+ voffcv = -0.10701 acde = 0.8 moin = 18.13
+ cgsl = {9.548271750000001E-12/sw_func_tox_lv_ratio} cgdl = {9.548271750000001E-12/sw_func_tox_lv_ratio} ijthsrev = 0.1
+ ijthsfwd = 0.1 xjbvs = 1 bvs = 12.69
+ jss = 2.1483E-5 jsws = 8.040000000000001E-10 cjs = {sw_psd_nw_cj}
+ mjs = 0.34629 mjsws = 0.29781 cjsws = {9.888891999999999E-11*sw_func_psd_nw_cj}
+ cjswgs = {2.39155046E-10*sw_func_psd_nw_cj} mjswgs = 0.9274 pbs = 0.6587
+ pbsws = 0.7418 pbswgs = 1.4338 xrcrg1 = 12
+ xrcrg2 = 1 rbpb = 50 rbpd = 50
+ rbps = 50 rbdb = 50 rbsb = 50
+ gbmin = 1E-12 tnom = 30 ute = -0.16467132300088
+ lute = -1.427567007550114E-7 kt1 = -0.45620503904216 lkt1 = -1.634479430716797E-8
+ kt1l = 0 kt2 = -0.040349144324356 lkt2 = -7.20772827667392E-9
+ ua1 = 1.4159172613352E-9 lua1 = 4.708289264257502E-16 ub1 = -8.959962135999941E-21
+ lub1 = -1.224117766644938E-24 uc1 = -2.1606649321236E-11 luc1 = 1.038808120716675E-17
+ at = 7.0857671813008E4 lat = 0.02052868205901 prt = 0
+ njs = 1.3632 xtis = 5.2 tpb = 2.0386E-3
+ tpbsw = 1.246E-3 tpbswg = 0 tcj = 1.2407E-3
+ tcjsw = 3.7357E-4 tcjswg = 2E-12 tvoff = 0
+ tvfbsdoff = 0 saref = 3E-6 sbref = 3E-6
+ wlod = 0 ku0 = 4.5E-8 kvsat = 0.5
+ kvth0 = 3.29E-8 tku0 = 0 llodku0 = 0
+ wlodku0 = 1 llodvth = 0 wlodvth = 1
+ lku0 = 0 wku0 = 2.5E-7 pku0 = 0
+ lkvth0 = 0 wkvth0 = 2E-7 pkvth0 = 0
+ stk2 = 0 lodk2 = 1 steta0 = 0
+ lodeta0 = 1

.model pshort_model.5 pmos
+ level = 54 lmin = 5E-7 lmax = 1E-6 wmin = 7E-6
+ wmax = 1.01E-3 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 4.23E-9
+ toxm = 4.23E-9 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 9.999999999999999E22 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {7.3039E-9+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {-1.3994E-8-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = -5.722E-9 dwb = -1.7864E-8 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = -1.0624270051384 lvth0 = 3.189929531261361E-8
+ k1 = 0.56285163226288 lk1 = -4.618105768145347E-8 k2 = -0.036139298542928
+ lk2 = 2.372902494638746E-8 k3 = -15.845 k3b = 2
+ w0 = 0 lpe0 = 0 lpeb = 0
+ vbm = -3 dvtp0 = 0 dvtp1 = 0
+ dvt0 = 4.4955 dvt1 = 0.294 dvt2 = 0.015
+ dvt0w = -4.9772 dvt1w = 1.1472E6 dvt2w = -8.96E-3
+ vfbsdoff = 0 u0 = 0.0102388475208 lu0 = -1.68615476841215E-9
+ ua = -6.448941519468001E-10 lua = -3.60086204608713E-16 ub = 1.00672124302384E-18
+ lub = 1.805592015719286E-25 uc = -5.9342542976688E-11 luc = 2.441319149781954E-17
+ ud = 0 up = 0 lp = 1
+ eu = 1.67 vsat = 5.97458806632E4 lvsat = 0.011826096628798
+ a0 = 0.99242407784 la0 = -4.351892401058587E-8 ags = 0.39408181584584
+ lags = 2.348729138113067E-7 b0 = 0 b1 = 0
+ keta = -0.0433129398494 lketa = 1.748385527110501E-8 a1 = 0
+ a2 = 1.0055976 la2 = -1.085530656288E-7 rdsw = 547.88
+ rdswmin = 0 rdw = 0 rdwmin = 0
+ rsw = 0 rswmin = 0 prwb = -0.32348
+ prwg = 0.1376 wr = 1 voff = -0.22937597595944
+ lvoff = -3.678114378007199E-9 voffl = 0 minv = 0
+ nfactor = 1.6385354519392 lnfactor = 2.608617009512568E-8 eta0 = 0.49
+ etab = -15.292603399365598 letab = 8.074278084374242E-6 dsub = 0.21844986818264
+ ldsub = 4.271303690666424E-8 cit = 1E-5 cdsc = 1.3E-4
+ cdscb = 7.8E-4 cdscd = 0 pclm = 0.61161503644472
+ lpclm = 6.066520638585094E-9 pdiblc1 = 0.723599095127128 lpdiblc1 = -3.61537833735426E-7
+ pdiblc2 = 4.3E-4 pdiblcb = 0.236063617142644 lpdiblcb = -2.434360570879102E-7
+ drout = 0.41525382127056 ldrout = 3.087389654149994E-7 pscbe1 = 8E8
+ pscbe2 = 8.713198730509598E-9 lpscbe2 = 2.285453447604983E-16 pvag = 0
+ delta = 0.01 fprout = 0 pdits = 0
+ pditsl = 0 pditsd = 0 lambda = 0
+ vtl = 0 lc = 5E-9 xn = 3
+ alpha0 = 9.1793747738312E-5 lalpha0 = -4.846594448205587E-11 alpha1 = -1.055976E-10
+ lalpha1 = 1.085530656288E-16 beta0 = 51.532746936979194 lbeta0 = -2.224334728221537E-5
+ aigbacc = 0.43 bigbacc = 0.054 cigbacc = 0.075
+ nigbacc = 1 aigbinv = 0.35 bigbinv = 0.03
+ cigbinv = 6E-3 eigbinv = 1.1 nigbinv = 3
+ aigc = 0.43 bigc = 0.054 cigc = 0.075
+ aigsd = 0.43 bigsd = 0.054 cigsd = 0.075
+ dlcig = 0 nigc = 1 poxedge = 1
+ pigcd = 1 ntox = 1 toxref = 4.23E-9
+ agidl = 1E-10 bgidl = 1.7182139032296E9 lbgidl = -370.63501159079
+ cgidl = 300 egidl = 0.1 noia = 1.5E42
+ noib = 0 noic = 0 em = 4.1E7
+ af = 1 ef = 1 kf = 0
+ lintnoi = -2E-7 tnoia = 2.5E7 tnoib = 0
+ ntnoi = 1 rnoia = 0.69 rnoib = 0.34
+ xpart = 0 cgso = {5.248925E-11/sw_func_tox_lv_ratio} cgdo = {5.248925E-11/sw_func_tox_lv_ratio}
+ cgbo = {0/sw_func_tox_lv_ratio} ckappas = 0.6 cf = 1.2E-11
+ clc = 1E-7 cle = 0.6 dlc = -3E-9
+ dwc = 0 vfbcv = -0.14469 noff = 3.9
+ voffcv = -0.10701 acde = 0.8 moin = 18.13
+ cgsl = {9.548271750000001E-12/sw_func_tox_lv_ratio} cgdl = {9.548271750000001E-12/sw_func_tox_lv_ratio} ijthsrev = 0.1
+ ijthsfwd = 0.1 xjbvs = 1 bvs = 12.69
+ jss = 2.1483E-5 jsws = 8.040000000000001E-10 cjs = {sw_psd_nw_cj}
+ mjs = 0.34629 mjsws = 0.29781 cjsws = {9.888891999999999E-11*sw_func_psd_nw_cj}
+ cjswgs = {2.39155046E-10*sw_func_psd_nw_cj} mjswgs = 0.9274 pbs = 0.6587
+ pbsws = 0.7418 pbswgs = 1.4338 xrcrg1 = 12
+ xrcrg2 = 1 rbpb = 50 rbpd = 50
+ rbps = 50 rbdb = 50 rbsb = 50
+ gbmin = 1E-12 tnom = 30 ute = -0.23309857548808
+ lute = -7.241430632519963E-8 kt1 = -0.43371464300408 lkt1 = -3.946465154956185E-8
+ kt1l = 0 kt2 = -0.03909512541676 lkt2 = -8.496844665455723E-9
+ ua1 = 3.3723123594224E-9 lua1 = -1.540321757666714E-15 ub1 = -2.9027539688824E-18
+ lub1 = 1.75066774676228E-24 uc1 = -4.9327926350544E-11 luc1 = 3.888522133797102E-17
+ at = 1.0754083678144E5 lat = -0.017181171330559 prt = 0
+ njs = 1.3632 xtis = 5.2 tpb = 2.0386E-3
+ tpbsw = 1.246E-3 tpbswg = 0 tcj = 1.2407E-3
+ tcjsw = 3.7357E-4 tcjswg = 2E-12 tvoff = 0
+ tvfbsdoff = 0 saref = 2.75E-6 sbref = 2.74E-6
+ wlod = 0 ku0 = 4.5E-8 kvsat = 0.5
+ kvth0 = 3.29E-8 tku0 = 0 llodku0 = 0
+ wlodku0 = 1 llodvth = 0 wlodvth = 1
+ lku0 = 0 wku0 = 2.5E-7 pku0 = 0
+ lkvth0 = 0 wkvth0 = 2E-7 pkvth0 = 0
+ stk2 = 0 lodk2 = 1 steta0 = 0
+ lodeta0 = 1

.model pshort_model.6 pmos
+ level = 54 lmin = 2.5E-7 lmax = 5E-7 wmin = 7E-6
+ wmax = 1.01E-3 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 4.23E-9
+ toxm = 4.23E-9 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 9.999999999999999E22 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {7.3039E-9+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {-1.3994E-8-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = -5.722E-9 dwb = -1.7864E-8 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = -1.0124385194416 lvth0 = 5.505974726531539E-9
+ k1 = 0.08709568447584 lk1 = 2.050123736787302E-7 k2 = 0.14027851671536
+ lk2 = -6.941746449620551E-8 k3 = -15.845 k3b = 2
+ w0 = 0 lpe0 = 0 lpeb = 0
+ vbm = -3 dvtp0 = 0 dvtp1 = 0
+ dvt0 = 4.4955 dvt1 = 0.294 dvt2 = 0.015
+ dvt0w = -4.9772 dvt1w = 1.1472E6 dvt2w = -8.96E-3
+ vfbsdoff = 0 u0 = 0.01008390899136 lu0 = -1.604349084130184E-9
+ ua = -5.189863622912E-10 lua = -4.265640066533939E-16 ub = 7.784653081887997E-19
+ lub = 3.01075596093612E-25 uc = -2.778294195410422E-11 luc = 7.750100873107581E-18
+ ud = 0 up = 0 lp = 1
+ eu = 1.67 vsat = 6.16513582256E4 lvsat = 0.010820027341582
+ a0 = 1.19308860166064 la0 = -1.49467384613598E-7 ags = -0.50603033730192
+ lags = 7.101213293274863E-7 b0 = 0 b1 = 0
+ keta = 0.069579111951392 lketa = -4.212179337509157E-8 a1 = 0
+ a2 = 0.8 rdsw = 547.88 rdswmin = 0
+ rdw = 0 rdwmin = 0 rsw = 0
+ rswmin = 0 prwb = -0.32348 prwg = 0.1376
+ wr = 1 voff = -0.20612908974192 lvoff = -1.595219133822314E-8
+ voffl = 0 minv = 0 nfactor = 1.3360896749344
+ lnfactor = 1.857739110043362E-7 eta0 = 1.032990803345882 leta0 = -2.866926282769854E-7
+ etab = 5.465032962355202E-3 letab = -2.918471073727998E-9 dsub = 0.1689577833808
+ ldsub = 6.88442637770182E-8 cit = 1E-5 cdsc = 1.3E-4
+ cdscb = 7.8E-4 cdscd = 0 pclm = 0.45686117965856
+ lpclm = 8.777469997539626E-8 pdiblc1 = -0.387531337591376 lpdiblc1 = 2.251257011747515E-7
+ pdiblc2 = -0.010312532689536 lpdiblc2 = 5.671928349682736E-9 pdiblcb = -0.3917928
+ lpdiblcb = 8.806459688640004E-8 drout = 1.59065746041392 ldrout = -3.118600512090249E-7
+ pscbe1 = 8E8 pscbe2 = 9.440251520520001E-9 lpscbe2 = -1.55329803731514E-16
+ pvag = 0 delta = 0.01 fprout = 0
+ pdits = 0 pditsl = 0 pditsd = 0
+ lambda = 0 vtl = 0 lc = 5E-9
+ xn = 3 alpha0 = -8.838017509640004E-9 lalpha0 = 4.719165988879806E-15
+ alpha1 = 2.111952E-10 lalpha1 = -5.870973125760002E-17 beta0 = 2.5236342748896
+ lbeta0 = 3.63287609401599E-6 aigbacc = 0.43 bigbacc = 0.054
+ cigbacc = 0.075 nigbacc = 1 aigbinv = 0.35
+ bigbinv = 0.03 cigbinv = 6E-3 eigbinv = 1.1
+ nigbinv = 3 aigc = 0.43 bigc = 0.054
+ cigc = 0.075 aigsd = 0.43 bigsd = 0.054
+ cigsd = 0.075 dlcig = 0 nigc = 1
+ poxedge = 1 pigcd = 1 ntox = 1
+ toxref = 4.23E-9 agidl = 1E-10 bgidl = 4.089569018911998E8
+ lbgidl = 320.63697403186916 cgidl = 560.2121596395841 lcgidl = -1.373888977437847E-4
+ egidl = 0.1 noia = 1.5E42 noib = 0
+ noic = 0 em = 4.1E7 af = 1
+ ef = 1 kf = 0 lintnoi = -2E-7
+ tnoia = 2.5E7 tnoib = 0 ntnoi = 1
+ rnoia = 0.69 rnoib = 0.34 xpart = 0
+ cgso = {5.248925E-11/sw_func_tox_lv_ratio} cgdo = {5.248925E-11/sw_func_tox_lv_ratio} cgbo = {0/sw_func_tox_lv_ratio}
+ ckappas = 0.6 cf = 1.2E-11 clc = 1E-7
+ cle = 0.6 dlc = -3E-9 dwc = 0
+ vfbcv = -0.14469 noff = 3.9 voffcv = -0.10701
+ acde = 0.8 moin = 18.13 cgsl = {9.548271750000001E-12/sw_func_tox_lv_ratio}
+ cgdl = {9.548271750000001E-12/sw_func_tox_lv_ratio} ijthsrev = 0.1 ijthsfwd = 0.1
+ xjbvs = 1 bvs = 12.69 jss = 2.1483E-5
+ jsws = 8.040000000000001E-10 cjs = {sw_psd_nw_cj} mjs = 0.34629
+ mjsws = 0.29781 cjsws = {9.888891999999999E-11*sw_func_psd_nw_cj} cjswgs = {2.39155046E-10*sw_func_psd_nw_cj}
+ mjswgs = 0.9274 pbs = 0.6587 pbsws = 0.7418
+ pbswgs = 1.4338 xrcrg1 = 12 xrcrg2 = 1
+ rbpb = 50 rbpd = 50 rbps = 50
+ rbdb = 50 rbsb = 50 gbmin = 1E-12
+ tnom = 30 ute = -0.378311652 lute = 4.256455516176021E-9
+ kt1 = -0.45237314112 lkt1 = -2.961318844633341E-8 kt1l = 0
+ kt2 = 0.019059258944 lkt2 = -3.920166175532468E-8 ua1 = 8.111838232E-10
+ lua1 = -1.880766240837216E-16 ub1 = 4.3553038656E-19 lub1 = -1.190633349904128E-26
+ uc1 = 9.125175919999995E-12 luc1 = 8.022684776351041E-18 at = 6.165657599999999E4
+ lat = 7.045167750912002E-3 prt = 0 njs = 1.3632
+ xtis = 5.2 tpb = 2.0386E-3 tpbsw = 1.246E-3
+ tpbswg = 0 tcj = 1.2407E-3 tcjsw = 3.7357E-4
+ tcjswg = 2E-12 tvoff = 0 tvfbsdoff = 0
+ saref = 1.75E-6 sbref = 1.74E-6 wlod = 0
+ ku0 = 4.5E-8 kvsat = 0.5 kvth0 = 3.29E-8
+ tku0 = 0 llodku0 = 0 wlodku0 = 1
+ llodvth = 0 wlodvth = 1 lku0 = 0
+ wku0 = 2.5E-7 pku0 = 0 lkvth0 = 0
+ wkvth0 = 2E-7 pkvth0 = 0 stk2 = 0
+ lodk2 = 1 steta0 = 0 lodeta0 = 1

.model pshort_model.7 pmos
+ level = 54 lmin = 1.8E-7 lmax = 2.5E-7 wmin = 7E-6
+ wmax = 1.01E-3 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 4.23E-9
+ toxm = 4.23E-9 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 9.999999999999999E22 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {7.3039E-9+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {-1.3994E-8-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = -5.722E-9 dwb = -1.7864E-8 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = -0.897340812171429 lvth0 = -2.648980672208888E-8
+ k1 = 0.237429301868572 lk1 = 1.632214320469595E-7 k2 = 0.109518224818628
+ lk2 = -6.08664724724169E-8 k3 = -15.845 k3b = 2
+ w0 = 0 lpe0 = 0 lpeb = 0
+ vbm = -3 dvtp0 = 0 dvtp1 = 0
+ dvt0 = 4.4955 dvt1 = 0.294 dvt2 = 0.015
+ dvt0w = -4.9772 dvt1w = 1.1472E6 dvt2w = -8.96E-3
+ vfbsdoff = 0 u0 = 6.034641789714285E-3 lu0 = -4.787013932790947E-10
+ ua = -1.399966414897142E-9 lua = -1.816621237895732E-16 ub = 1.256083153794286E-18
+ lub = 1.68303566429434E-25 uc = -7.826224615577139E-14 luc = 4.853237045440658E-20
+ ud = 0 up = 0 lp = 1
+ eu = 1.67 vsat = 1.329054374742857E5 lvsat = -8.987751640601732E-3
+ a0 = 1.023500970640572 la0 = -1.023240582415912E-7 ags = 4.42094239888
+ lags = -6.595179676582535E-7 b0 = 0 b1 = 0
+ keta = -0.255963735087943 lketa = 4.837521158767906E-8 a1 = 0
+ a2 = 0.884075316078286 la2 = -2.337192896597052E-8 rdsw = 547.88
+ rdswmin = 0 rdw = 0 rdwmin = 0
+ rsw = 0 rswmin = 0 prwb = -0.32348
+ prwg = 0.1376 wr = 1 voff = -0.067040389644
+ lvoff = -5.461718090104376E-8 voffl = 0 minv = 0
+ nfactor = 1.685791809142858 lnfactor = 8.856091411999532E-8 eta0 = -0.500893996689577
+ leta0 = 1.397089395152718E-7 etab = 0.150037252567531 letab = -4.310781325733173E-8
+ dsub = 0.813536297068 ldsub = -1.103408280858592E-7 cit = 1E-5
+ cdsc = 1.3E-4 cdscb = 7.8E-4 cdscd = 0
+ pclm = 1.177407606724571 lpclm = -1.125285601918301E-7 pdiblc1 = 1.122642611480571
+ lpdiblc1 = -1.946845345798611E-7 pdiblc2 = 0.027672729654789 lpdiblc2 = -4.887518758891365E-9
+ pdiblcb = -0.075 drout = -0.960132607944571 ldrout = 3.972289783138154E-7
+ pscbe1 = 7.9999646E8 pscbe2 = 7.932893943971429E-9 lpscbe2 = 2.636975142580706E-16
+ pvag = 0 delta = 0.01 fprout = 0
+ pdits = 0 pditsl = 0 pditsd = 0
+ lambda = 0 vtl = 0 lc = 5E-9
+ xn = 3 alpha0 = 3.202149110585715E-8 lalpha0 = -6.639287092125016E-15
+ alpha1 = -2.971257142857143E-10 lalpha1 = 8.259738306285714E-17 beta0 = 36.351762977919996
+ lbeta0 = -5.770937747882025E-6 aigbacc = 0.43 bigbacc = 0.054
+ cigbacc = 0.075 nigbacc = 1 aigbinv = 0.35
+ bigbinv = 0.03 cigbinv = 6E-3 eigbinv = 1.1
+ nigbinv = 3 aigc = 0.43 bigc = 0.054
+ cigc = 0.075 aigsd = 0.43 bigsd = 0.054
+ cigsd = 0.075 dlcig = 0 nigc = 1
+ poxedge = 1 pigcd = 1 ntox = 1
+ toxref = 4.23E-9 agidl = 6.135698839028571E-11 lagidl = 1.074229351136126E-17
+ bgidl = 3.233344075354285E9 lbgidl = -464.50876754478713 cgidl = -629.3291415699427
+ lcgidl = 1.932893094968493E-4 egidl = 0.1 noia = 1.5E42
+ noib = 0 noic = 0 em = 4.1E7
+ af = 1 ef = 1 kf = 0
+ lintnoi = -2E-7 tnoia = 2.5E7 tnoib = 0
+ ntnoi = 1 rnoia = 0.69 rnoib = 0.34
+ xpart = 0 cgso = {5.248925E-11/sw_func_tox_lv_ratio} cgdo = {5.248925E-11/sw_func_tox_lv_ratio}
+ cgbo = {0/sw_func_tox_lv_ratio} ckappas = 0.6 cf = 1.2E-11
+ clc = 1E-7 cle = 0.6 dlc = -3E-9
+ dwc = 0 vfbcv = -0.14469 noff = 3.9
+ voffcv = -0.10701 acde = 0.8 moin = 18.13
+ cgsl = {9.548271750000001E-12/sw_func_tox_lv_ratio} cgdl = {9.548271750000001E-12/sw_func_tox_lv_ratio} ijthsrev = 0.1
+ ijthsfwd = 0.1 xjbvs = 1 bvs = 12.69
+ jss = 2.1483E-5 jsws = 8.040000000000001E-10 cjs = {sw_psd_nw_cj}
+ mjs = 0.34629 mjsws = 0.29781 cjsws = {9.888891999999999E-11*sw_func_psd_nw_cj}
+ cjswgs = {2.39155046E-10*sw_func_psd_nw_cj} mjswgs = 0.9274 pbs = 0.6587
+ pbsws = 0.7418 pbswgs = 1.4338 xrcrg1 = 12
+ xrcrg2 = 1 rbpb = 50 rbpd = 50
+ rbps = 50 rbdb = 50 rbsb = 50
+ gbmin = 1E-12 tnom = 30 ute = -0.5501892
+ lute = 5.20363513296E-8 kt1 = -0.5589 kt1l = 0
+ kt2 = -0.12196 ua1 = 1.3462E-10 ub1 = 3.927E-19
+ uc1 = 3.7985E-11 at = 2.325916E5 lat = -0.0404727177008
+ prt = 0 njs = 1.3632 xtis = 5.2
+ tpb = 2.0386E-3 tpbsw = 1.246E-3 tpbswg = 0
+ tcj = 1.2407E-3 tcjsw = 3.7357E-4 tcjswg = 2E-12
+ tvoff = 0 tvfbsdoff = 0 saref = 1.25E-6
+ sbref = 1.24E-6 wlod = 0 ku0 = 4.5E-8
+ kvsat = 0.5 kvth0 = 3.29E-8 tku0 = 0
+ llodku0 = 0 wlodku0 = 1 llodvth = 0
+ wlodvth = 1 lku0 = 0 wku0 = 2.5E-7
+ pku0 = 0 lkvth0 = 0 wkvth0 = 2E-7
+ pkvth0 = 0 stk2 = 0 lodk2 = 1
+ steta0 = 0 lodeta0 = 1

.model pshort_model.8 pmos
+ level = 54 lmin = 1.5E-7 lmax = 1.8E-7 wmin = 7E-6
+ wmax = 1.01E-3 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 4.23E-9
+ toxm = 4.23E-9 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 9.999999999999999E22 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {7.3039E-9+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {-1.3994E-8-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = -5.722E-9 dwb = -1.7864E-8 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = -0.8585156044 lvth0 = -3.456498403605279E-8
+ k1 = -0.556924842106666 lk1 = 3.284375617440813E-7 k2 = 0.480439082930666
+ lk2 = -1.380135599094234E-7 k3 = -15.845 k3b = 2
+ w0 = 0 lpe0 = 0 lpeb = 0
+ vbm = -3 dvtp0 = 0 dvtp1 = 0
+ dvt0 = 4.4955 dvt1 = 0.294 dvt2 = 0.015
+ dvt0w = -4.9772 dvt1w = 1.1472E6 dvt2w = -8.96E-3
+ vfbsdoff = 0 u0 = 6.933818203999995E-3 lu0 = -6.657192973335512E-10
+ ua = -8.685443885733356E-10 lua = -2.921915282006091E-16 ub = 7.070587317599995E-19
+ lub = 2.824940579195012E-25 uc = 2.975755702373331E-13 luc = -2.963738530156245E-20
+ ud = 0 up = 0 lp = 1
+ eu = 1.67 vsat = 2.769247034266666E5 lvsat = -0.038942030727506
+ a0 = -1.110903038712 la0 = 3.416063628556314E-7 ags = 1.25
+ b0 = 0 b1 = 0 keta = -0.108048302823173
+ lketa = 1.761057666179416E-8 a1 = 0 a2 = -0.579795937515999
+ la2 = 2.810957253265977E-7 rdsw = 547.88 rdswmin = 0
+ rdw = 0 rdwmin = 0 rsw = 0
+ rswmin = 0 prwb = -0.32348 prwg = 0.1376
+ wr = 1 voff = 0.036059445901333 lvoff = -7.606070949644647E-8
+ voffl = 0 minv = 0 nfactor = -0.020528251999997
+ lnfactor = 4.434550109969754E-7 eta0 = -0.807748139174666 leta0 = 2.035309189024604E-7
+ etab = -0.292823200157333 letab = 4.900184658400741E-8 dsub = 0.419602642290666
+ ldsub = -2.840735509603115E-8 cit = 1E-5 cdsc = 1.3E-4
+ cdscb = 7.8E-4 cdscd = 0 pclm = 2.476238444478666
+ lpclm = -3.826697884746287E-7 pdiblc1 = 1.178029696558666 lpdiblc1 = -2.062043836310838E-7
+ pdiblc2 = 0.026384736551627 lpdiblc2 = -4.619631649350925E-9 pdiblcb = -0.501673309421253
+ lpdiblcb = 8.874292827990758E-8 drout = 0.651497248421334 ldrout = 6.20293077479837E-8
+ pscbe1 = 8.835736127773333E8 lpscbe1 = -17.382308574331994 pscbe2 = 1.035851282288E-8
+ lpscbe2 = -2.408021051283657E-16 pvag = 0 delta = 0.01
+ fprout = 0 pdits = 0 pditsl = 0
+ pditsd = 0 lambda = 0 vtl = 0
+ lc = 5E-9 xn = 3 alpha0 = 1E-10
+ alpha1 = 1E-10 beta0 = 15.8918131392 lbeta0 = -1.515513700826329E-6
+ aigbacc = 0.43 bigbacc = 0.054 cigbacc = 0.075
+ nigbacc = 1 aigbinv = 0.35 bigbinv = 0.03
+ cigbinv = 6E-3 eigbinv = 1.1 nigbinv = 3
+ aigc = 0.43 bigc = 0.054 cigc = 0.075
+ aigsd = 0.43 bigsd = 0.054 cigsd = 0.075
+ dlcig = 0 nigc = 1 poxedge = 1
+ pigcd = 1 ntox = 1 toxref = 4.23E-9
+ agidl = 1.901670270893333E-10 lagidl = -1.604864881757625E-17 bgidl = 7.280064512133335E8
+ lbgidl = 56.571394225041196 cgidl = 300 egidl = 0.1
+ noia = 1.5E42 noib = 0 noic = 0
+ em = 4.1E7 af = 1 ef = 1
+ kf = 0 lintnoi = -2E-7 tnoia = 2.5E7
+ tnoib = 0 ntnoi = 1 rnoia = 0.69
+ rnoib = 0.34 xpart = 0 cgso = {5.248925E-11/sw_func_tox_lv_ratio}
+ cgdo = {5.248925E-11/sw_func_tox_lv_ratio} cgbo = {0/sw_func_tox_lv_ratio} ckappas = 0.6
+ cf = 1.2E-11 clc = 1E-7 cle = 0.6
+ dlc = -3E-9 dwc = 0 vfbcv = -0.14469
+ noff = 3.9 voffcv = -0.10701 acde = 0.8
+ moin = 18.13 cgsl = {9.548271750000001E-12/sw_func_tox_lv_ratio} cgdl = {9.548271750000001E-12/sw_func_tox_lv_ratio}
+ ijthsrev = 0.1 ijthsfwd = 0.1 xjbvs = 1
+ bvs = 12.69 jss = 2.1483E-5 jsws = 8.040000000000001E-10
+ cjs = {sw_psd_nw_cj} mjs = 0.34629 mjsws = 0.29781
+ cjsws = {9.888891999999999E-11*sw_func_psd_nw_cj} cjswgs = {2.39155046E-10*sw_func_psd_nw_cj} mjswgs = 0.9274
+ pbs = 0.6587 pbsws = 0.7418 pbswgs = 1.4338
+ xrcrg1 = 12 xrcrg2 = 1 rbpb = 50
+ rbpd = 50 rbps = 50 rbdb = 50
+ rbsb = 50 gbmin = 1E-12 tnom = 30
+ ute = -0.3 kt1 = 0.21890756 lkt1 = -1.617746387892799E-7
+ kt1l = 0 kt2 = -0.12196 ua1 = 1.3462E-10
+ ub1 = 3.927E-19 uc1 = 3.7985E-11 at = 3.8E4
+ prt = 0 njs = 1.3632 xtis = 5.2
+ tpb = 2.0386E-3 tpbsw = 1.246E-3 tpbswg = 0
+ tcj = 1.2407E-3 tcjsw = 3.7357E-4 tcjswg = 2E-12
+ tvoff = 0 tvfbsdoff = 0 saref = 1.1E-6
+ sbref = 1.1E-6 wlod = 0 ku0 = 4.5E-8
+ kvsat = 0.5 kvth0 = 3.29E-8 tku0 = 0
+ llodku0 = 0 wlodku0 = 1 llodvth = 0
+ wlodvth = 1 lku0 = 0 wku0 = 2.5E-7
+ pku0 = 0 lkvth0 = 0 wkvth0 = 2E-7
+ pkvth0 = 0 stk2 = 0 lodk2 = 1
+ steta0 = 0 lodeta0 = 1

.model pshort_model.9 pmos
+ level = 54 lmin = 8E-6 lmax = 2.02E-5 wmin = 5E-6
+ wmax = 7E-6 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 4.23E-9
+ toxm = 4.23E-9 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 9.999999999999999E22 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {7.3039E-9+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {-1.3994E-8-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = -5.722E-9 dwb = -1.7864E-8 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = -1.070814813024892 wvth0 = 7.866461831191605E-8
+ k1 = 0.444261859177239 wk1 = -6.829149357931748E-8 k2 = 0.015623434959989
+ wk2 = 2.901669777838879E-8 k3 = -15.845 k3b = 2
+ w0 = 0 lpe0 = 0 lpeb = 0
+ vbm = -3 dvtp0 = 0 dvtp1 = 0
+ dvt0 = 4.4955 dvt1 = 0.294 dvt2 = 0.015
+ dvt0w = -4.9772 dvt1w = 1.1472E6 dvt2w = -8.96E-3
+ vfbsdoff = 0 u0 = 0.01077223375746 wu0 = -2.065117743417805E-9
+ ua = -5.908449854809399E-10 wua = 1.745668754204094E-16 ub = 9.43061924020675E-19
+ wub = -7.011562287780338E-26 uc = -7.483094472841781E-11 wuc = 5.784589818864008E-17
+ ud = 0 up = 0 lp = 1
+ eu = 1.67 vsat = 1.603125E5 a0 = 1.3425676466503
+ wa0 = -7.386887860793633E-7 ags = 0.221790026409061 wags = 3.028009363091169E-8
+ b0 = 0 b1 = 0 keta = 0.03003246861336
+ wketa = -1.739604290434864E-7 a1 = 0 a2 = 1.223159949392132
+ wa2 = -1.562352465936194E-6 rdsw = 547.88 rdswmin = 0
+ rdw = 0 rdwmin = 0 rsw = 0
+ rswmin = 0 prwb = -0.32348 prwg = 0.1376
+ wr = 1 voff = -0.269379060845788 wvoff = 8.603635733260264E-8
+ voffl = 0 minv = 0 nfactor = 0.77913338195144
+ wnfactor = 3.901602923444549E-6 eta0 = 0.08 etab = -0.07
+ dsub = 0.56 cit = 1E-5 cdsc = 1.3E-4
+ cdscb = 7.8E-4 cdscd = 0 pclm = -0.561230562720794
+ wpclm = 3.931052954664842E-6 pdiblc1 = 0.39 pdiblc2 = 9.92920113806031E-3
+ wpdiblc2 = -4.865992589279954E-8 pdiblcb = -0.025 drout = 0.56
+ pscbe1 = 8E8 pscbe2 = 1.012148770893988E-8 wpscbe2 = -5.206861812043943E-15
+ pvag = 0 delta = 0.01 fprout = 0
+ pdits = 0 pditsl = 0 pditsd = 0
+ lambda = 0 vtl = 0 lc = 5E-9
+ xn = 3 alpha0 = 1E-10 alpha1 = 1E-10
+ beta0 = 0.396943770666869 wbeta0 = 2.968412258986038E-5 aigbacc = 0.43
+ bigbacc = 0.054 cigbacc = 0.075 nigbacc = 1
+ aigbinv = 0.35 bigbinv = 0.03 cigbinv = 6E-3
+ eigbinv = 1.1 nigbinv = 3 aigc = 0.43
+ bigc = 0.054 cigc = 0.075 aigsd = 0.43
+ bigsd = 0.054 cigsd = 0.075 dlcig = 0
+ nigc = 1 poxedge = 1 pigcd = 1
+ ntox = 1 toxref = 4.23E-9 agidl = 1E-10
+ bgidl = 2.804225407656603E8 wbgidl = 6.291459561391775E3 cgidl = 300
+ egidl = 0.1 noia = 1.5E42 noib = 0
+ noic = 0 em = 4.1E7 af = 1
+ ef = 1 kf = 0 lintnoi = -2E-7
+ tnoia = 2.5E7 tnoib = 0 ntnoi = 1
+ rnoia = 0.69 rnoib = 0.34 xpart = 0
+ cgso = {5.248925E-11/sw_func_tox_lv_ratio} cgdo = {5.248925E-11/sw_func_tox_lv_ratio} cgbo = {0/sw_func_tox_lv_ratio}
+ ckappas = 0.6 cf = 1.2E-11 clc = 1E-7
+ cle = 0.6 dlc = -3E-9 dwc = 0
+ vfbcv = -0.14469 noff = 3.9 voffcv = -0.10701
+ acde = 0.8 moin = 18.13 cgsl = {9.548271750000001E-12/sw_func_tox_lv_ratio}
+ cgdl = {9.548271750000001E-12/sw_func_tox_lv_ratio} ijthsrev = 0.1 ijthsfwd = 0.1
+ xjbvs = 1 bvs = 12.69 jss = 2.1483E-5
+ jsws = 8.040000000000001E-10 cjs = {sw_psd_nw_cj} mjs = 0.34629
+ mjsws = 0.29781 cjsws = {9.888891999999999E-11*sw_func_psd_nw_cj} cjswgs = {2.39155046E-10*sw_func_psd_nw_cj}
+ mjswgs = 0.9274 pbs = 0.6587 pbsws = 0.7418
+ pbswgs = 1.4338 xrcrg1 = 12 xrcrg2 = 1
+ rbpb = 50 rbpd = 50 rbps = 50
+ rbdb = 50 rbsb = 50 gbmin = 1E-12
+ tnom = 30 ute = -0.775332799574229 wute = 3.044183622961982E-6
+ kt1 = -0.479524993031196 wkt1 = 2.167217443251707E-7 kt1l = 0
+ kt2 = 0.099528252454443 wkt2 = -7.481274885642141E-7 ua1 = 7.405564963019101E-10
+ wua1 = 6.076198025953308E-15 ub1 = -8.348099522392428E-20 wub1 = -3.334958992094562E-24
+ uc1 = -6.582460621904258E-10 wuc1 = 3.839633023429716E-15 at = 9.314342649E4
+ wat = -0.015671213904519 prt = 0 njs = 1.3632
+ xtis = 5.2 tpb = 2.0386E-3 tpbsw = 1.246E-3
+ tpbswg = 0 tcj = 1.2407E-3 tcjsw = 3.7357E-4
+ tcjswg = 2E-12 tvoff = 0 tvfbsdoff = 0
+ saref = 3E-6 sbref = 3E-6 wlod = 0
+ ku0 = 4.5E-8 kvsat = 0.5 kvth0 = 3.29E-8
+ tku0 = 0 llodku0 = 0 wlodku0 = 1
+ llodvth = 0 wlodvth = 1 lku0 = 0
+ wku0 = 2.5E-7 pku0 = 0 lkvth0 = 0
+ wkvth0 = 2E-7 pkvth0 = 0 stk2 = 0
+ lodk2 = 1 steta0 = 0 lodeta0 = 1

.model pshort_model.10 pmos
+ level = 54 lmin = 4E-6 lmax = 8E-6 wmin = 5E-6
+ wmax = 7E-6 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 4.23E-9
+ toxm = 4.23E-9 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 9.999999999999999E22 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {7.3039E-9+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {-1.3994E-8-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = -5.722E-9 dwb = -1.7864E-8 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = -1.072176032955128 lvth0 = 1.092785726529274E-8
+ wvth0 = 6.314027965773959E-8 pvth0 = 1.246292044236647E-13 k1 = 0.417770816632546
+ lk1 = 2.126697716562863E-7 wk1 = 1.422413822506808E-7 pk1 = -1.690155400768717E-12
+ k2 = 0.023858077730997 lk2 = -6.610761334994251E-8 wk2 = -3.739241008545311E-8
+ pk2 = 5.331315210216283E-13 k3 = -15.845 k3b = 2
+ w0 = 0 lpe0 = 0 lpeb = 0
+ vbm = -3 dvtp0 = 0 dvtp1 = 0
+ dvt0 = 4.4955 dvt1 = 0.294 dvt2 = 0.015
+ dvt0w = -4.9772 dvt1w = 1.1472E6 dvt2w = -8.96E-3
+ vfbsdoff = 0 u0 = 0.011988142905293 lu0 = -9.761304047894323E-9
+ wu0 = -1.18825694443716E-8 pu0 = 7.881438444583668E-14 ua = -2.35694865293704E-10
+ lua = -2.851140903061689E-15 wua = -2.386602524851971E-15 pua = 2.056103721135386E-20
+ ub = 6.956340199309337E-19 lub = 1.986348244897594E-24 wub = 1.623271880129644E-24
+ pub = -1.359449455349375E-29 uc = -9.304491999719303E-11 luc = 1.462215748900243E-16
+ wuc = 1.384471240505861E-16 puc = -6.470656740049924E-22 ud = 0
+ up = 0 lp = 1 eu = 1.67
+ vsat = 2.762846165846647E5 lvsat = -0.93102276027629 wvsat = -0.058323220384757
+ pvsat = 4.682181133701822E-7 a0 = 1.622216337228062 la0 = -2.245016332173988E-6
+ wa0 = -2.049254587980394E-6 pa0 = 1.052120653087185E-11 ags = 0.179857368541926
+ lags = 3.366348741654659E-7 wags = -1.820686337764218E-7 pags = 1.704733035441345E-12
+ b0 = 0 b1 = 0 keta = 0.073052536666315
+ lketa = -3.453645900883041E-7 wketa = -3.604162754817509E-7 pketa = 1.49686529773623E-12
+ a1 = 0 a2 = 1.649280748950161 la2 = -3.420892665402261E-6
+ wa2 = -3.135636712076543E-6 pa2 = 1.263030704860377E-11 rdsw = 547.88
+ rdswmin = 0 rdw = 0 rdwmin = 0
+ rsw = 0 rswmin = 0 prwb = -0.32348
+ prwg = 0.1376 wr = 1 voff = -0.300303243065369
+ lvoff = 2.482589637686089E-7 wvoff = 2.32599566539057E-7 pvoff = -1.176607684750905E-12
+ voffl = 0 minv = 0 nfactor = 0.220392379615384
+ lnfactor = 4.485566061861827E-6 wnfactor = 6.726342759344261E-6 pnfactor = -2.267697750572486E-11
+ eta0 = 0.08 etab = -0.07 dsub = 0.56
+ cit = 1E-5 cdsc = 1.3E-4 cdscb = 7.8E-4
+ cdscd = 0 pclm = -1.546484603803385 lpclm = 7.909607618762542E-6
+ wpclm = 7.77393072983995E-6 ppclm = -3.085057666457246E-11 pdiblc1 = 0.39
+ pdiblc2 = 0.019645712020002 lpdiblc2 = -7.800403276209932E-8 wpdiblc2 = -9.679330227408829E-8
+ ppdiblc2 = 3.864141679884695E-13 pdiblcb = -0.025 drout = 0.56
+ pscbe1 = 8E8 pscbe2 = 1.377023184625808E-8 lpscbe2 = -2.929207414946093E-14
+ wpscbe2 = -2.534656528941901E-14 ppscbe2 = 1.616812978399253E-19 pvag = 0
+ delta = 0.01 fprout = 0 pdits = 0
+ pditsl = 0 pditsd = 0 lambda = 0
+ vtl = 0 lc = 5E-9 xn = 3
+ alpha0 = 1E-10 alpha1 = 1E-10 beta0 = -3.699146609143646
+ lbeta0 = 3.288336441603427E-5 wbeta0 = 4.850391097930663E-5 pbeta0 = -1.510850353530138E-10
+ aigbacc = 0.43 bigbacc = 0.054 cigbacc = 0.075
+ nigbacc = 1 aigbinv = 0.35 bigbinv = 0.03
+ cigbinv = 6E-3 eigbinv = 1.1 nigbinv = 3
+ aigc = 0.43 bigc = 0.054 cigc = 0.075
+ aigsd = 0.43 bigsd = 0.054 cigsd = 0.075
+ dlcig = 0 nigc = 1 poxedge = 1
+ pigcd = 1 ntox = 1 toxref = 4.23E-9
+ agidl = 4.504973268132962E-11 lagidl = 4.411400866310781E-16 wagidl = 2.739486340784143E-16
+ pagidl = -2.199256346997901E-21 bgidl = 7.773279455744288E8 lbgidl = -3.989150626939935E3
+ wbgidl = 4.094159919609314E3 pbgidl = 0.017639895156634 cgidl = 300
+ egidl = 0.1 noia = 1.5E42 noib = 0
+ noic = 0 em = 4.1E7 af = 1
+ ef = 1 kf = 0 lintnoi = -2E-7
+ tnoia = 2.5E7 tnoib = 0 ntnoi = 1
+ rnoia = 0.69 rnoib = 0.34 xpart = 0
+ cgso = {5.248925E-11/sw_func_tox_lv_ratio} cgdo = {5.248925E-11/sw_func_tox_lv_ratio} cgbo = {0/sw_func_tox_lv_ratio}
+ ckappas = 0.6 cf = 1.2E-11 clc = 1E-7
+ cle = 0.6 dlc = -3E-9 dwc = 0
+ vfbcv = -0.14469 noff = 3.9 voffcv = -0.10701
+ acde = 0.8 moin = 18.13 cgsl = {9.548271750000001E-12/sw_func_tox_lv_ratio}
+ cgdl = {9.548271750000001E-12/sw_func_tox_lv_ratio} ijthsrev = 0.1 ijthsfwd = 0.1
+ xjbvs = 1 bvs = 12.69 jss = 2.1483E-5
+ jsws = 8.040000000000001E-10 cjs = {sw_psd_nw_cj} mjs = 0.34629
+ mjsws = 0.29781 cjsws = {9.888891999999999E-11*sw_func_psd_nw_cj} cjswgs = {2.39155046E-10*sw_func_psd_nw_cj}
+ mjswgs = 0.9274 pbs = 0.6587 pbsws = 0.7418
+ pbswgs = 1.4338 xrcrg1 = 12 xrcrg2 = 1
+ rbpb = 50 rbpd = 50 rbps = 50
+ rbdb = 50 rbsb = 50 gbmin = 1E-12
+ tnom = 30 ute = -1.349052455176396 lute = 4.605814510538336E-6
+ wute = 6.109625141083179E-6 pute = -2.460932772217875E-11 kt1 = -0.487713346053629
+ lkt1 = 6.573599980385881E-8 wkt1 = 3.92157800188842E-7 pkt1 = -1.408398551240883E-12
+ kt1l = 0 kt2 = 0.157972924743657 lkt2 = -4.691931278017501E-7
+ wkt2 = -1.035019342953909E-6 pkt2 = 2.303164364338221E-12 ua1 = -5.226090295054814E-11
+ lua1 = 6.364728567389943E-15 wua1 = 8.91427444653555E-15 pua1 = -2.278404344751719E-20
+ ub1 = 4.0123251243327E-19 lub1 = -3.891274222909864E-24 wub1 = -4.894166706308628E-24
+ pub1 = 1.251730081921795E-29 uc1 = -1.195561529593474E-9 luc1 = 4.313562124526062E-15
+ wuc1 = 7.734635182845605E-15 puc1 = -3.126903059576484E-20 at = 9.337414290628923E4
+ lat = -1.852188621372986E-3 wat = -0.038517698755876 pat = 1.834113062288736E-7
+ prt = 0 njs = 1.3632 xtis = 5.2
+ tpb = 2.0386E-3 tpbsw = 1.246E-3 tpbswg = 0
+ tcj = 1.2407E-3 tcjsw = 3.7357E-4 tcjswg = 2E-12
+ tvoff = 0 tvfbsdoff = 0 saref = 3E-6
+ sbref = 3E-6 wlod = 0 ku0 = 4.5E-8
+ kvsat = 0.5 kvth0 = 3.29E-8 tku0 = 0
+ llodku0 = 0 wlodku0 = 1 llodvth = 0
+ wlodvth = 1 lku0 = 0 wku0 = 2.5E-7
+ pku0 = 0 lkvth0 = 0 wkvth0 = 2E-7
+ pkvth0 = 0 stk2 = 0 lodk2 = 1
+ steta0 = 0 lodeta0 = 1

.model pshort_model.11 pmos
+ level = 54 lmin = 2E-6 lmax = 4E-6 wmin = 5E-6
+ wmax = 7E-6 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 4.23E-9
+ toxm = 4.23E-9 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 9.999999999999999E22 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {7.3039E-9+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {-1.3994E-8-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = -5.722E-9 dwb = -1.7864E-8 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = -1.07803369344703 lvth0 = 3.452244343475155E-8
+ wvth0 = 9.348943101665388E-8 pvth0 = 2.383186939774301E-15 k1 = 0.515778983259006
+ lk1 = -1.82105947417098E-7 wk1 = -6.392108224254744E-7 pk1 = 1.457524702240381E-12
+ k2 = -8.710277499466772E-3 lk2 = 6.507733069810342E-8 wk2 = 2.235984216695884E-7
+ pk2 = -5.181364173976979E-13 k3 = -15.845 k3b = 2
+ w0 = 0 lpe0 = 0 lpeb = 0
+ vbm = -3 dvtp0 = 0 dvtp1 = 0
+ dvt0 = 4.4955 dvt1 = 0.294 dvt2 = 0.015
+ dvt0w = -4.9772 dvt1w = 1.1472E6 dvt2w = -8.96E-3
+ vfbsdoff = 0 u0 = 8.459350659924987E-3 lu0 = 4.452628770941498E-9
+ wu0 = 2.589465088637918E-8 pu0 = -7.335180571978349E-14 ua = -1.296687962484564E-9
+ lua = 1.422526560505929E-15 wua = 7.444229534666704E-15 pua = -1.903743635440264E-20
+ ub = 1.415787157137852E-18 lub = -9.144199499342259E-25 wub = -4.631517636063488E-24
+ pub = 1.159972256025799E-29 uc = -6.229406098266247E-11 luc = 2.235748378980339E-17
+ wuc = -1.299118672128172E-16 puc = 4.338811224961011E-22 ud = 0
+ up = 0 lp = 1 eu = 1.67
+ vsat = 3.673887558067053E4 lvsat = 0.033864609938907 wvsat = 0.116646440769514
+ pvsat = -2.365575821232844E-7 a0 = 1.097480235062625 la0 = -1.313856094848319E-7
+ wa0 = 5.180830391014298E-7 pa0 = 1.800013770377899E-13 ags = -0.070590837458984
+ lags = 1.34543724255866E-6 wags = 1.152627209053603E-6 pags = -3.671405803127883E-12
+ b0 = 0 b1 = 0 keta = -8.989592400778765E-3
+ lketa = -1.489987871159874E-8 wketa = 2.462232333177754E-8 pketa = -5.406555782147676E-14
+ a1 = 0 a2 = 0.8 rdsw = 547.88
+ rdswmin = 0 rdw = 0 rdwmin = 0
+ rsw = 0 rswmin = 0 prwb = -0.32348
+ prwg = 0.1376 wr = 1 voff = -0.254605045408927
+ lvoff = 6.418717198683341E-8 wvoff = 3.505193409987713E-9 pvoff = -2.538182989194935E-13
+ voffl = 0 minv = 0 nfactor = 0.928009366123205
+ lnfactor = 1.635293331612165E-6 wnfactor = 4.095202257642372E-6 pnfactor = -1.207877513855567E-11
+ eta0 = 0.160612527827676 leta0 = -3.247062947395438E-7 peta0 = 1.358366776413661E-19
+ etab = -0.140472582538707 letab = 2.838627167949205E-7 petab = 7.111868507750544E-22
+ dsub = 0.8641982 ldsub = -1.2253066992216E-6 cit = 1E-5
+ cdsc = 1.3E-4 cdscb = 7.8E-4 cdscd = 0
+ pclm = 1.028039343348187 lpclm = -2.460543946076622E-6 wpclm = -3.935761274253052E-6
+ ppclm = 1.63159222116101E-11 pdiblc1 = 0.39 pdiblc2 = 4.71776621692122E-4
+ lpdiblc2 = -7.71651064930894E-10 wpdiblc2 = -3.446350211975349E-9 ppdiblc2 = 1.041376524570332E-14
+ pdiblcb = -0.025 drout = 0.56 pscbe1 = 7.723676175051484E8
+ lpscbe1 = 111.30290510067232 wpscbe1 = 196.14053409842074 ppscbe1 = -7.900517176620296E-4
+ pscbe2 = 5.321470778700365E-9 lpscbe2 = 4.739434045528769E-15 wpscbe2 = 2.071143048888577E-14
+ ppscbe2 = -2.383975645913702E-20 pvag = 0 delta = 0.01
+ fprout = 0 pdits = 0 pditsl = 0
+ pditsd = 0 lambda = 0 vtl = 0
+ lc = 5E-9 xn = 3 alpha0 = 1E-10
+ alpha1 = 1E-10 beta0 = 0.927342922078164 lbeta0 = 1.424792010214719E-5
+ wbeta0 = 2.07302233985774E-5 pbeta0 = -3.921295506208746E-11 aigbacc = 0.43
+ bigbacc = 0.054 cigbacc = 0.075 nigbacc = 1
+ aigbinv = 0.35 bigbinv = 0.03 cigbinv = 6E-3
+ eigbinv = 1.1 nigbinv = 3 aigc = 0.43
+ bigc = 0.054 cigc = 0.075 aigsd = 0.43
+ bigsd = 0.054 cigsd = 0.075 dlcig = 0
+ nigc = 1 poxedge = 1 pigcd = 1
+ ntox = 1 toxref = 4.23E-9 agidl = 2.099005346373408E-10
+ lagidl = -2.228769654381114E-16 wagidl = -5.478972681568286E-16 pagidl = 1.11112908505483E-21
+ bgidl = -8.594637480716248E8 lbgidl = 2.603826673566044E3 wbgidl = 1.241105920082468E4
+ pbgidl = -0.01586047534531 cgidl = 300 egidl = 0.1
+ noia = 1.5E42 noib = 0 noic = 0
+ em = 4.1E7 af = 1 ef = 1
+ kf = 0 lintnoi = -2E-7 tnoia = 2.5E7
+ tnoib = 0 ntnoi = 1 rnoia = 0.69
+ rnoib = 0.34 xpart = 0 cgso = {5.248925E-11/sw_func_tox_lv_ratio}
+ cgdo = {5.248925E-11/sw_func_tox_lv_ratio} cgbo = {0/sw_func_tox_lv_ratio} ckappas = 0.6
+ cf = 1.2E-11 clc = 1E-7 cle = 0.6
+ dlc = -3E-9 dwc = 0 vfbcv = -0.14469
+ noff = 3.9 voffcv = -0.10701 acde = 0.8
+ moin = 18.13 cgsl = {9.548271750000001E-12/sw_func_tox_lv_ratio} cgdl = {9.548271750000001E-12/sw_func_tox_lv_ratio}
+ ijthsrev = 0.1 ijthsfwd = 0.1 xjbvs = 1
+ bvs = 12.69 jss = 2.1483E-5 jsws = 8.040000000000001E-10
+ cjs = {sw_psd_nw_cj} mjs = 0.34629 mjsws = 0.29781
+ cjsws = {9.888891999999999E-11*sw_func_psd_nw_cj} cjswgs = {2.39155046E-10*sw_func_psd_nw_cj} mjswgs = 0.9274
+ pbs = 0.6587 pbsws = 0.7418 pbswgs = 1.4338
+ xrcrg1 = 12 xrcrg2 = 1 rbpb = 50
+ rbpd = 50 rbps = 50 rbdb = 50
+ rbsb = 50 gbmin = 1E-12 tnom = 30
+ ute = -0.326588997179382 lute = 4.873439712878543E-7 wute = 1.05394818483942E-6
+ pute = -4.245121610552365E-12 kt1 = -0.481217021021369 lkt1 = 3.956888052981599E-8
+ wkt1 = 1.037301404862631E-7 pkt1 = -2.466153990908117E-13 kt1l = 0
+ kt2 = 0.125810850004869 lkt2 = -3.39644676698805E-7 wkt2 = -9.171063352940923E-7
+ pkt2 = 1.82821218444057E-12 ua1 = 1.030333228276962E-9 lua1 = 2.00405239793511E-15
+ wua1 = 9.185209249293568E-15 pua1 = -2.387536558180885E-20 ub1 = -3.551467258727138E-19
+ lub1 = -8.445877275642207E-25 wub1 = -4.724680198682162E-24 pub1 = 1.183461120033663E-29
+ uc1 = 9.563768158812432E-11 luc1 = -8.873728037228821E-16 wuc1 = -2.362153701442745E-15
+ puc1 = 9.40071386868202E-21 at = 1.013841037720225E5 lat = -0.034116214869016
+ wat = 0.039496388202415 pat = -1.308284998700779E-7 prt = 0
+ njs = 1.3632 xtis = 5.2 tpb = 2.0386E-3
+ tpbsw = 1.246E-3 tpbswg = 0 tcj = 1.2407E-3
+ tcjsw = 3.7357E-4 tcjswg = 2E-12 tvoff = 0
+ tvfbsdoff = 0 saref = 3E-6 sbref = 3E-6
+ wlod = 0 ku0 = 4.5E-8 kvsat = 0.5
+ kvth0 = 3.29E-8 tku0 = 0 llodku0 = 0
+ wlodku0 = 1 llodvth = 0 wlodvth = 1
+ lku0 = 0 wku0 = 2.5E-7 pku0 = 0
+ lkvth0 = 0 wkvth0 = 2E-7 pkvth0 = 0
+ stk2 = 0 lodk2 = 1 steta0 = 0
+ lodeta0 = 1

.model pshort_model.12 pmos
+ level = 54 lmin = 1E-6 lmax = 2E-6 wmin = 5E-6
+ wmax = 7E-6 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 4.23E-9
+ toxm = 4.23E-9 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 9.999999999999999E22 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {7.3039E-9+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {-1.3994E-8-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = -5.722E-9 dwb = -1.7864E-8 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = -1.084032632112787 lvth0 = 4.668821906164124E-8
+ wvth0 = 1.401372309255739E-7 pvth0 = -9.221799150191655E-14 k1 = 0.324438550909221
+ lk1 = 2.059301533030792E-7 wk1 = 2.102881690677843E-7 pk1 = -2.652490585200498E-13
+ k2 = 0.066384155545189 lk2 = -8.721327838326241E-8 wk2 = -1.034463962339315E-7
+ pk2 = 1.451065487728256E-13 k3 = -15.845 k3b = 2
+ w0 = 0 lpe0 = 0 lpeb = 0
+ vbm = -3 dvtp0 = 0 dvtp1 = 0
+ dvt0 = 4.4955 dvt1 = 0.294 dvt2 = 0.015
+ dvt0w = -4.9772 dvt1w = 1.1472E6 dvt2w = -8.96E-3
+ vfbsdoff = 0 u0 = 0.011047114778513 lu0 = -7.953258083856701E-10
+ wu0 = -8.810888958004278E-9 pu0 = -2.969387381851981E-15 ua = -5.350455367405788E-10
+ lua = -1.220751391937637E-16 wua = -1.489215698699699E-15 pua = -9.205166224783767E-22
+ ub = 9.290061085013814E-19 lub = 7.276617532795277E-26 wub = 8.960192482805799E-25
+ pub = 3.899440892508332E-31 uc = -5.362968853891524E-11 luc = 4.786240446353324E-18
+ wuc = 7.434289670444955E-17 puc = 1.96549123290511E-23 ud = 0
+ up = 0 lp = 1 eu = 1.67
+ vsat = -7.579273164358202E4 lvsat = 0.262077359010405 wvsat = 0.774814082332604
+ pvsat = -1.571313661201533E-6 a0 = 0.463295678794674 la0 = 1.154733060411897E-6
+ wa0 = 5.801309848539633E-6 pa0 = -1.053431919378117E-11 ags = 1.946855431203339
+ lags = -2.745919580933307E-6 wags = -1.100558524137924E-5 pags = 2.098530314780052E-11
+ b0 = 0 b1 = 0 keta = -0.072443434075034
+ lketa = 1.137837507576898E-7 wketa = 4.593776099694486E-7 pketa = -9.35744062059234E-13
+ a1 = 0 a2 = 0.44095503215532 la2 = 7.281388862493966E-7
+ wa2 = 1.789979982142118E-6 pa2 = -3.630057924024429E-12 rdsw = 547.88
+ rdswmin = 0 rdw = 0 rdwmin = 0
+ rsw = 0 rswmin = 0 prwb = -0.32348
+ prwg = 0.1376 wr = 1 voff = -0.208292079609894
+ lvoff = -2.973496689801676E-8 wvoff = -2.773258053589153E-7 pvoff = 3.157035966118575E-13
+ voffl = 0 minv = 0 nfactor = 2.065514468729105
+ lnfactor = -6.715533664113694E-7 wnfactor = -5.580946532134427E-6 pnfactor = 7.544338493326201E-12
+ eta0 = -0.502700135655351 leta0 = 1.020483827052073E-6 peta0 = -6.933410634732136E-20
+ etab = 26.70210614008915 letab = -5.415256482174971E-5 wetab = -1.331191203419064E-4
+ petab = 2.699639786242951E-10 dsub = 0.26 cit = 1E-5
+ cdsc = 1.3E-4 cdscb = 7.8E-4 cdscd = 0
+ pclm = -1.51475066928458 lpclm = 2.696203686062479E-6 wpclm = 1.185669062005024E-5
+ ppclm = -1.571098072061425E-11 pdiblc1 = 0.432576358597428 lpdiblc1 = -8.634434431928156E-8
+ wpdiblc1 = -1.674705271292171E-7 ppdiblc1 = 3.396282193717268E-13 pdiblc2 = -2.569285774587309E-4
+ lpdiblc2 = 7.061543344846458E-10 wpdiblc2 = 3.424608372019852E-9 ppdiblc2 = -3.520456311135944E-15
+ pdiblcb = -0.049980264489432 lpdiblcb = 5.065967662139373E-8 wpdiblcb = 3.217186511283275E-10
+ ppdiblcb = -6.524415638644346E-16 drout = 0.6468349600767 ldrout = -1.761002570160257E-7
+ wdrout = -1.723831271902054E-6 pdrout = 3.495909133442104E-12 pscbe1 = 8.552647649897032E8
+ lpscbe1 = -56.81151523223502 wpscbe1 = -392.2810681968415 ppscbe1 = 4.032602307335347E-4
+ pscbe2 = 1.923792875317121E-9 lpscbe2 = 1.162988406145515E-14 wpscbe2 = 4.905155843707296E-14
+ ppscbe2 = -8.131319585652528E-20 pvag = 0 delta = 0.01
+ fprout = 0 pdits = 0 pditsl = 0
+ pditsd = 0 lambda = 0 vtl = 0
+ lc = 5E-9 xn = 3 alpha0 = -1.60303557730188E-4
+ lalpha0 = 3.250938942329286E-10 walpha0 = 7.991766048795493E-10 palpha0 = -1.620720564576467E-15
+ alpha1 = 4.590449678446798E-10 lalpha1 = -7.281388862493967E-16 walpha1 = -1.789979982142118E-15
+ palpha1 = 3.63005792402443E-21 beta0 = -68.32365600446198 lbeta0 = 1.546881149131835E-4
+ wbeta0 = 3.780865783801057E-4 pbeta0 = -7.639273546883671E-10 aigbacc = 0.43
+ bigbacc = 0.054 cigbacc = 0.075 nigbacc = 1
+ aigbinv = 0.35 bigbinv = 0.03 cigbinv = 6E-3
+ eigbinv = 1.1 nigbinv = 3 aigc = 0.43
+ bigc = 0.054 cigc = 0.075 aigsd = 0.43
+ bigsd = 0.054 cigsd = 0.075 dlcig = 0
+ nigc = 1 poxedge = 1 pigcd = 1
+ ntox = 1 toxref = 4.23E-9 agidl = 1E-10
+ bgidl = -9.81367553268815E8 lbgidl = 2.851046127660285E3 wbgidl = 1.242828733741204E4
+ pbgidl = -0.015895413799572 cgidl = 300 egidl = 0.1
+ noia = 1.5E42 noib = 0 noic = 0
+ em = 4.1E7 af = 1 ef = 1
+ kf = 0 lintnoi = -2E-7 tnoia = 2.5E7
+ tnoib = 0 ntnoi = 1 rnoia = 0.69
+ rnoib = 0.34 xpart = 0 cgso = {5.248925E-11/sw_func_tox_lv_ratio}
+ cgdo = {5.248925E-11/sw_func_tox_lv_ratio} cgbo = {0/sw_func_tox_lv_ratio} ckappas = 0.6
+ cf = 1.2E-11 clc = 1E-7 cle = 0.6
+ dlc = -3E-9 dwc = 0 vfbcv = -0.14469
+ noff = 3.9 voffcv = -0.10701 acde = 0.8
+ moin = 18.13 cgsl = {9.548271750000001E-12/sw_func_tox_lv_ratio} cgdl = {9.548271750000001E-12/sw_func_tox_lv_ratio}
+ ijthsrev = 0.1 ijthsfwd = 0.1 xjbvs = 1
+ bvs = 12.69 jss = 2.1483E-5 jsws = 8.040000000000001E-10
+ cjs = {sw_psd_nw_cj} mjs = 0.34629 mjsws = 0.29781
+ cjsws = {9.888891999999999E-11*sw_func_psd_nw_cj} cjswgs = {2.39155046E-10*sw_func_psd_nw_cj} mjswgs = 0.9274
+ pbs = 0.6587 pbsws = 0.7418 pbswgs = 1.4338
+ xrcrg1 = 12 xrcrg2 = 1 rbpb = 50
+ rbpd = 50 rbps = 50 rbdb = 50
+ rbsb = 50 gbmin = 1E-12 tnom = 30
+ ute = 0.300064203004743 lute = -7.835011988471481E-7 wute = -3.246359918422578E-6
+ pute = 4.475851619165728E-12 kt1 = -0.455903412914567 lkt1 = -1.176681294748212E-8
+ wkt1 = -2.106976799005254E-9 pkt1 = -3.197899528169492E-14 kt1l = 0
+ kt2 = -0.036716377258421 lkt2 = -1.004141013558113E-8 wkt2 = -2.537630272680005E-8
+ pkt2 = 1.979437915449192E-14 ua1 = 2.246181378111194E-9 lua1 = -4.616730597509175E-16
+ wua1 = -5.799720485266921E-15 pua1 = 6.513892100723003E-21 ub1 = -4.277360238529569E-19
+ lub1 = -6.973775023318636E-25 wub1 = 2.92531503506435E-24 pub1 = -3.679487333758487E-30
+ uc1 = -6.807951057229347E-10 luc1 = 6.872235717504977E-16 wuc1 = 4.604689901678467E-15
+ puc1 = -4.727961356324558E-21 at = -8.949404975502074E4 lat = 0.352982389945985
+ wat = 1.12011966509788 pat = -2.322319537934759E-6 prt = 0
+ njs = 1.3632 xtis = 5.2 tpb = 2.0386E-3
+ tpbsw = 1.246E-3 tpbswg = 0 tcj = 1.2407E-3
+ tcjsw = 3.7357E-4 tcjswg = 2E-12 tvoff = 0
+ tvfbsdoff = 0 saref = 3E-6 sbref = 3E-6
+ wlod = 0 ku0 = 4.5E-8 kvsat = 0.5
+ kvth0 = 3.29E-8 tku0 = 0 llodku0 = 0
+ wlodku0 = 1 llodvth = 0 wlodvth = 1
+ lku0 = 0 wku0 = 2.5E-7 pku0 = 0
+ lkvth0 = 0 wkvth0 = 2E-7 pkvth0 = 0
+ stk2 = 0 lodk2 = 1 steta0 = 0
+ lodeta0 = 1

.model pshort_model.13 pmos
+ level = 54 lmin = 5E-7 lmax = 1E-6 wmin = 5E-6
+ wmax = 7E-6 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 4.23E-9
+ toxm = 4.23E-9 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 9.999999999999999E22 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {7.3039E-9+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {-1.3994E-8-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = -5.722E-9 dwb = -1.7864E-8 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = -1.065934911151001 lvth0 = 2.808397908557691E-8
+ wvth0 = 2.450409929875314E-8 pvth0 = 2.665148021287564E-14 k1 = 0.592920162830969
+ lk1 = -7.006572197313452E-8 wk1 = -2.100404788957883E-7 pk1 = 1.668437476427273E-13
+ k2 = -0.05439092955334 lk2 = 3.694205979700415E-8 wk2 = 1.274948008974081E-7
+ pk2 = -9.229823058382593E-14 k3 = -15.845 k3b = 2
+ w0 = 0 lpe0 = 0 lpeb = 0
+ vbm = -3 dvtp0 = 0 dvtp1 = 0
+ dvt0 = 4.4955 dvt1 = 0.294 dvt2 = 0.015
+ dvt0w = -4.9772 dvt1w = 1.1472E6 dvt2w = -8.96E-3
+ vfbsdoff = 0 u0 = 0.013044231637226 lu0 = -2.848337973740075E-9
+ wu0 = -1.959670832488469E-8 pu0 = 8.11830549746868E-15 ua = -3.552447620872214E-11
+ lua = -6.355767951677859E-16 wua = -4.256686179817298E-15 pua = 1.924409822464742E-21
+ ub = 7.177820785419627E-19 lub = 2.899019434378754E-25 wub = 2.018353385846224E-24
+ pub = -7.63801936156998E-31 uc = -8.367664269366062E-11 luc = 3.567414875398173E-17
+ wuc = 1.699832303569628E-16 puc = -7.866220298172874E-23 ud = 0
+ up = 0 lp = 1 eu = 1.67
+ vsat = 2.796377393938912E5 lvsat = -0.103300900050465 wvsat = -1.536030874820872
+ pvsat = 8.042072246127552E-7 a0 = 2.28083725199641 la0 = -7.136778663406088E-7
+ wa0 = -9.000071337129426E-6 pa0 = 4.681323048512392E-12 ags = -2.250038573770686
+ lags = 1.56843709345193E-6 wags = 1.847021794548824E-5 pags = -9.31546881866101E-12
+ b0 = 0 b1 = 0 keta = 0.079484376266709
+ lketa = -4.239621513989763E-8 wketa = -8.57787414178404E-7 pketa = 4.182857767844686E-13
+ a1 = 0 a2 = 1.524753840146547 la2 = -3.859932827798884E-7
+ wa2 = -3.626509950501015E-6 pa2 = 1.93802872885352E-12 rdsw = 547.88
+ rdswmin = 0 rdw = 0 rdwmin = 0
+ rsw = 0 rswmin = 0 prwb = -0.32348
+ prwg = 0.1376 wr = 1 voff = -0.244832686193965
+ lvoff = 7.828338183129591E-9 wvoff = 1.079711831099117E-7 pvoff = -8.037708397023495E-14
+ voffl = 0 minv = 0 nfactor = 1.040035020201209
+ lnfactor = 3.82627200921925E-7 wnfactor = 4.180760247559194E-6 pnfactor = -2.490578935717484E-12
+ eta0 = 0.49 etab = -53.406092014421716 letab = 2.81977015827096E-5
+ wetab = 2.662376660864018E-4 petab = -1.405700055425685E-10 dsub = 0.199057618246563
+ ldsub = 6.264803713395194E-8 wdsub = 1.354624714439213E-7 pdsub = -1.392537950946938E-13
+ cit = 1E-5 cdsc = 1.3E-4 cdscb = 7.8E-4
+ cdscd = 0 pclm = 1.622117103152611 lpclm = -5.284587415896848E-7
+ wpclm = -7.058753254865183E-6 ppclm = 3.733868597472311E-12 pdiblc1 = 0.624709378761775
+ lpdiblc1 = -2.838547834519881E-7 wpdiblc1 = 6.907834533587474E-7 ppdiblc1 = -5.426465735221348E-13
+ pdiblc2 = 4.3E-4 pdiblcb = 0.236155728978863 lpdiblcb = -2.434846910320922E-7
+ wpdiblcb = -6.434373022566939E-10 ppdiblcb = 3.397271743439072E-16 drout = -0.078299360153399
+ ldrout = 5.693291225686727E-7 wdrout = 3.447662543804109E-6 pdrout = -1.820324451178044E-12
+ pscbe1 = 8E8 pscbe2 = -3.885259444036076E-9 lpscbe2 = 1.76015201371224E-14
+ wpscbe2 = 8.800517146449761E-14 ppscbe2 = -1.213570426053615E-19 pvag = 0
+ delta = 0.01 fprout = 0 pdits = 0
+ pditsl = 0 pditsd = 0 lambda = 0
+ vtl = 0 lc = 5E-9 xn = 3
+ alpha0 = 3.206074154603761E-4 lalpha0 = -1.69276815275293E-10 walpha0 = -1.598353209759098E-9
+ palpha0 = 8.439113145142867E-16 alpha1 = -6.1808993568936E-10 lalpha1 = 3.791428689647537E-16
+ walpha1 = 3.579959964284236E-15 palpha1 = -1.890175901622505E-21 beta0 = 158.99900912053818
+ lbeta0 = -7.899685696333516E-5 wbeta0 = -7.506939896201879E-4 pbeta0 = 3.964455238491186E-10
+ aigbacc = 0.43 bigbacc = 0.054 cigbacc = 0.075
+ nigbacc = 1 aigbinv = 0.35 bigbinv = 0.03
+ cigbinv = 6E-3 eigbinv = 1.1 nigbinv = 3
+ aigc = 0.43 bigc = 0.054 cigc = 0.075
+ aigsd = 0.43 bigsd = 0.054 cigsd = 0.075
+ dlcig = 0 nigc = 1 poxedge = 1
+ pigcd = 1 ntox = 1 toxref = 4.23E-9
+ agidl = 1E-10 bgidl = 3.146032936686658E9 lbgidl = -1.391872047208063E3
+ wbgidl = -9.973875939322475E3 pbgidl = 7.13374122295202E-3 cgidl = 300
+ egidl = 0.1 noia = 1.5E42 noib = 0
+ noic = 0 em = 4.1E7 af = 1
+ ef = 1 kf = 0 lintnoi = -2E-7
+ tnoia = 2.5E7 tnoib = 0 ntnoi = 1
+ rnoia = 0.69 rnoib = 0.34 xpart = 0
+ cgso = {5.248925E-11/sw_func_tox_lv_ratio} cgdo = {5.248925E-11/sw_func_tox_lv_ratio} cgbo = {0/sw_func_tox_lv_ratio}
+ ckappas = 0.6 cf = 1.2E-11 clc = 1E-7
+ cle = 0.6 dlc = -3E-9 dwc = 0
+ vfbcv = -0.14469 noff = 3.9 voffcv = -0.10701
+ acde = 0.8 moin = 18.13 cgsl = {9.548271750000001E-12/sw_func_tox_lv_ratio}
+ cgdl = {9.548271750000001E-12/sw_func_tox_lv_ratio} ijthsrev = 0.1 ijthsfwd = 0.1
+ xjbvs = 1 bvs = 12.69 jss = 2.1483E-5
+ jsws = 8.040000000000001E-10 cjs = {sw_psd_nw_cj} mjs = 0.34629
+ mjsws = 0.29781 cjsws = {9.888891999999999E-11*sw_func_psd_nw_cj} cjswgs = {2.39155046E-10*sw_func_psd_nw_cj}
+ mjswgs = 0.9274 pbs = 0.6587 pbsws = 0.7418
+ pbswgs = 1.4338 xrcrg1 = 12 xrcrg2 = 1
+ rbpb = 50 rbpd = 50 rbps = 50
+ rbdb = 50 rbsb = 50 gbmin = 1E-12
+ tnom = 30 ute = -0.420594685599675 lute = -4.267250926846928E-8
+ wute = 1.309733865103879E-6 pute = -2.077581171740672E-13 kt1 = -0.423938544205404
+ lkt1 = -4.462631440207726E-8 wkt1 = -6.828988429470145E-8 pkt1 = 3.605623942899083E-14
+ kt1l = 0 kt2 = -0.037293607233421 lkt2 = -9.448024648040302E-9
+ wkt2 = -1.258431106605161E-8 pkt2 = 6.644365231142455E-15 ua1 = 3.187989212252771E-9
+ lua1 = -1.429840211554448E-15 wua1 = 1.287569474518179E-15 pua1 = -7.717569304565617E-22
+ ub1 = -2.620271122607641E-18 lub1 = 1.556522268766767E-24 wub1 = -1.973253471001496E-24
+ pub1 = 1.35618230765513E-30 uc1 = -5.093259110282094E-11 luc1 = 3.973246507119622E-17
+ wuc1 = 1.120921264417033E-17 puc1 = -5.918329765570204E-24 at = 4.319241851544403E5
+ lat = -0.183029298522122 wat = -2.265944911534639 pat = 1.158514214068551E-6
+ prt = 0 njs = 1.3632 xtis = 5.2
+ tpb = 2.0386E-3 tpbsw = 1.246E-3 tpbswg = 0
+ tcj = 1.2407E-3 tcjsw = 3.7357E-4 tcjswg = 2E-12
+ tvoff = 0 tvfbsdoff = 0 saref = 2.75E-6
+ sbref = 2.74E-6 wlod = 0 ku0 = 4.5E-8
+ kvsat = 0.5 kvth0 = 3.29E-8 tku0 = 0
+ llodku0 = 0 wlodku0 = 1 llodvth = 0
+ wlodvth = 1 lku0 = 0 wku0 = 2.5E-7
+ pku0 = 0 lkvth0 = 0 wkvth0 = 2E-7
+ pkvth0 = 0 stk2 = 0 lodk2 = 1
+ steta0 = 0 lodeta0 = 1

.model pshort_model.14 pmos
+ level = 54 lmin = 2.5E-7 lmax = 5E-7 wmin = 5E-6
+ wmax = 7E-6 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 4.23E-9
+ toxm = 4.23E-9 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 9.999999999999999E22 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {7.3039E-9+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {-1.3994E-8-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = -5.722E-9 dwb = -1.7864E-8 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = -1.041034332957549 lvth0 = 1.493677260637241E-8
+ wvth0 = 1.997529726869592E-7 pvth0 = -6.58778219496165E-14 k1 = 0.051491016399681
+ lk1 = 2.158023701928279E-7 wk1 = 2.487125706627861E-7 pk1 = -7.537235748760526E-14
+ k2 = 0.159319176640184 lk2 = -7.58943117519023E-8 wk2 = -1.330064773217213E-7
+ pk2 = 4.524331830053575E-14 k3 = -15.845 k3b = 2
+ w0 = 0 lpe0 = 0 lpeb = 0
+ vbm = -3 dvtp0 = 0 dvtp1 = 0
+ dvt0 = 4.4955 dvt1 = 0.294 dvt2 = 0.015
+ dvt0w = -4.9772 dvt1w = 1.1472E6 dvt2w = -8.96E-3
+ vfbsdoff = 0 u0 = 0.011384237934039 lu0 = -1.971881218381624E-9
+ wu0 = -9.083307653620744E-9 pu0 = 2.567356103849362E-15 ua = -3.145111580591476E-10
+ lua = -4.882751749909435E-16 wua = -1.428339496735986E-15 pua = 4.310767139580061E-22
+ ub = 6.557725272402706E-19 lub = 3.226422424105532E-25 wub = 8.57057195034164E-25
+ pub = -1.506514829625202E-31 uc = -3.406880545732416E-11 luc = 9.481805987242905E-18
+ wuc = 4.390922188565717E-17 puc = -1.209663939698099E-23 ud = 0
+ up = 0 lp = 1 eu = 1.67
+ vsat = 1.994317573907722E4 lvsat = 0.033814713224512 wvsat = 0.291348012617533
+ pvsat = -1.606268994080735E-7 a0 = 1.270529017630105 la0 = -1.802472422940124E-7
+ wa0 = -5.409516776778551E-7 pa0 = 2.150093777578765E-13 ags = -0.161307728479942
+ lags = 4.656122719085609E-7 wags = -2.4080226228287E-6 pags = 1.707991662523514E-12
+ b0 = 0 b1 = 0 keta = 0.036472868525052
+ lketa = -1.968665519039556E-8 wketa = 2.31260094601656E-7 pketa = -1.567182392812977E-13
+ a1 = 0 a2 = 0.786672191085626 la2 = 3.704970944489045E-9
+ wa2 = 9.309997243355974E-8 pa2 = -2.588067513686041E-14 rdsw = 547.88
+ rdswmin = 0 rdw = 0 rdwmin = 0
+ rsw = 0 rswmin = 0 prwb = -0.32348
+ prwg = 0.1376 wr = 1 voff = -0.198053973684804
+ lvoff = -1.687026067715739E-8 wvoff = -5.640785271947362E-8 pvoff = 6.413074399250521E-15
+ voffl = 0 minv = 0 nfactor = 1.51612745620061
+ lnfactor = 1.312561078234732E-7 wnfactor = -1.257634512962296E-6 pnfactor = 3.808282371007358E-13
+ eta0 = 2.195850754915217 leta0 = -9.006687283861753E-7 weta0 = -8.12303283538481E-6
+ peta0 = 4.288863860689155E-12 etab = 0.015331155178636 letab = -8.168793761346463E-9
+ wetab = -6.891873317385243E-8 petab = 3.667556314957306E-14 dsub = 0.22030846578562
+ ldsub = 5.142784464350054E-8 wdsub = -3.587046563353064E-7 pdsub = 1.216605183672051E-13
+ cit = 1E-5 cdsc = 1.3E-4 cdscb = 7.8E-4
+ cdscd = 0 pclm = 0.228955171086373 lpclm = 2.071140405981044E-7
+ wpclm = 1.59201285461329E-6 ppclm = -8.336320991390086E-13 pdiblc1 = -0.436001593357445
+ lpdiblc1 = 2.761878812952948E-7 wpdiblc1 = 3.385837465603033E-7 ppdiblc1 = -3.566893547290381E-13
+ pdiblc2 = -0.019973891339189 lpdiblc2 = 1.077300978039594E-8 wpdiblc2 = 6.748837935269147E-8
+ ppdiblc2 = -3.563305443766886E-14 pdiblcb = -0.25320487931064 lpdiblcb = 1.489183781746625E-8
+ wpdiblcb = -9.680909801976738E-7 ppdiblcb = 5.111404204526093E-13 drout = 2.364847974238716
+ ldrout = -7.206233522223514E-7 wdrout = -5.408024376585724E-6 pdrout = 2.855371974544743E-12
+ pscbe1 = 8E8 pscbe2 = 6.575235951027063E-8 lpscbe2 = -1.916630701932408E-14
+ wpscbe2 = -3.933621599171617E-13 ppscbe2 = 1.32799131956178E-19 pvag = 0
+ delta = 0.01 fprout = 0 pdits = 0
+ pditsl = 0 pditsd = 0 lambda = 0
+ vtl = 0 lc = 5E-9 xn = 3
+ alpha0 = -7.80495931169916E-9 lalpha0 = 4.173723657065415E-15 walpha0 = -7.21631667804204E-15
+ palpha0 = 3.81012861020606E-21 alpha1 = 2.111952E-10 lalpha1 = -5.870973125760002E-17
+ beta0 = 2.53564170559846 lbeta0 = 3.613923471344025E-6 wbeta0 = -8.387661281571656E-8
+ pbeta0 = 1.323915025822886E-13 aigbacc = 0.43 bigbacc = 0.054
+ cigbacc = 0.075 nigbacc = 1 aigbinv = 0.35
+ bigbinv = 0.03 cigbinv = 6E-3 eigbinv = 1.1
+ nigbinv = 3 aigc = 0.43 bigc = 0.054
+ cigc = 0.075 aigsd = 0.43 bigsd = 0.054
+ cigsd = 0.075 dlcig = 0 nigc = 1
+ poxedge = 1 pigcd = 1 ntox = 1
+ toxref = 4.23E-9 agidl = 1E-10 bgidl = -9.908631051759352E7
+ lbgidl = 321.5119738848155 wbgidl = 3.548881093223328E3 pbgidl = -6.112217147772304E-6
+ cgidl = 485.5250392742439 lcgidl = -9.795499443632947E-5 wcgidl = 5.217188280405083E-4
+ pcgidl = -2.754612805794519E-10 egidl = 0.1 noia = 1.5E42
+ noib = 0 noic = 0 em = 4.1E7
+ af = 1 ef = 1 kf = 0
+ lintnoi = -2E-7 tnoia = 2.5E7 tnoib = 0
+ ntnoi = 1 rnoia = 0.69 rnoib = 0.34
+ xpart = 0 cgso = {5.248925E-11/sw_func_tox_lv_ratio} cgdo = {5.248925E-11/sw_func_tox_lv_ratio}
+ cgbo = {0/sw_func_tox_lv_ratio} ckappas = 0.6 cf = 1.2E-11
+ clc = 1E-7 cle = 0.6 dlc = -3E-9
+ dwc = 0 vfbcv = -0.14469 noff = 3.9
+ voffcv = -0.10701 acde = 0.8 moin = 18.13
+ cgsl = {9.548271750000001E-12/sw_func_tox_lv_ratio} cgdl = {9.548271750000001E-12/sw_func_tox_lv_ratio} ijthsrev = 0.1
+ ijthsfwd = 0.1 xjbvs = 1 bvs = 12.69
+ jss = 2.1483E-5 jsws = 8.040000000000001E-10 cjs = {sw_psd_nw_cj}
+ mjs = 0.34629 mjsws = 0.29781 cjsws = {9.888891999999999E-11*sw_func_psd_nw_cj}
+ cjswgs = {2.39155046E-10*sw_func_psd_nw_cj} mjswgs = 0.9274 pbs = 0.6587
+ pbsws = 0.7418 pbswgs = 1.4338 xrcrg1 = 12
+ xrcrg2 = 1 rbpb = 50 rbpd = 50
+ rbps = 50 rbdb = 50 rbsb = 50
+ gbmin = 1E-12 tnom = 30 ute = -0.480706468446889
+ lute = -1.093420926653464E-8 wute = 7.152679521285289E-7 pute = 1.061127512859617E-13
+ kt1 = -0.477596142685464 lkt1 = -1.629574629578746E-8 wkt1 = 1.761925583959766E-7
+ pkt1 = -9.302755652237489E-14 kt1l = 0 kt2 = 0.029203894738461
+ lkt2 = -4.455790771917062E-8 wkt2 = -7.086425975046967E-8 pkt2 = 3.741547877713098E-14
+ ua1 = 9.57125756545949E-10 lua1 = -2.519710773027146E-16 wua1 = -1.019461642847712E-15
+ pua1 = 4.463278151392184E-22 ub1 = 2.990830114142123E-19 lub1 = 1.51383182528367E-26
+ wub1 = 9.531384300538588E-25 pub1 = -1.889174993992847E-31 uc1 = -5.432591768841658E-11
+ luc1 = 4.152410078847169E-17 wuc1 = 4.43230774373703E-16 puc1 = -2.340205301000227E-22
+ at = 8.50865142454885E3 lat = 0.040529022300856 wat = 0.371259097775545
+ pat = -2.338978563991141E-7 prt = 0 njs = 1.3632
+ xtis = 5.2 tpb = 2.0386E-3 tpbsw = 1.246E-3
+ tpbswg = 0 tcj = 1.2407E-3 tcjsw = 3.7357E-4
+ tcjswg = 2E-12 tvoff = 0 tvfbsdoff = 0
+ saref = 1.75E-6 sbref = 1.74E-6 wlod = 0
+ ku0 = 4.5E-8 kvsat = 0.5 kvth0 = 3.29E-8
+ tku0 = 0 llodku0 = 0 wlodku0 = 1
+ llodvth = 0 wlodvth = 1 lku0 = 0
+ wku0 = 2.5E-7 pku0 = 0 lkvth0 = 0
+ wkvth0 = 2E-7 pkvth0 = 0 stk2 = 0
+ lodk2 = 1 steta0 = 0 lodeta0 = 1

.model pshort_model.15 pmos
+ level = 54 lmin = 1.8E-7 lmax = 2.5E-7 wmin = 5E-6
+ wmax = 7E-6 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 4.23E-9
+ toxm = 4.23E-9 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 9.999999999999999E22 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {7.3039E-9+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {-1.3994E-8-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = -5.722E-9 dwb = -1.7864E-8 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = -0.843499238756393 lvth0 = -3.997561316041861E-8
+ wvth0 = -3.761045069691203E-7 pvth0 = 9.420364710501829E-14 k1 = 0.345431055681784
+ lk1 = 1.340905665528748E-7 wk1 = -7.544346086731341E-7 pk1 = 2.034905206016286E-13
+ k2 = 0.069870084609664 lk2 = -5.102853755652208E-8 wk2 = 2.769578093602044E-7
+ pk2 = -6.872183382559942E-14 k3 = -15.845 k3b = 2
+ w0 = 0 lpe0 = 0 lpeb = 0
+ vbm = -3 dvtp0 = 0 dvtp1 = 0
+ dvt0 = 4.4955 dvt1 = 0.294 dvt2 = 0.015
+ dvt0w = -4.9772 dvt1w = 1.1472E6 dvt2w = -8.96E-3
+ vfbsdoff = 0 u0 = 4.765536881480205E-3 lu0 = -1.319617501830446E-10
+ wu0 = 8.865195526960053E-9 pu0 = -2.422112398313932E-15 ua = -1.431358861916722E-9
+ lua = -1.778049154909841E-16 wua = 2.192885545494858E-16 pua = -2.694411276273975E-23
+ ub = 9.027273581772006E-19 lub = 2.539917628680579E-25 wub = 2.468328818528385E-24
+ pub = -5.985656590344318E-31 uc = 1.739813078361896E-13 luc = -3.727782003048978E-20
+ wuc = -1.762020154555723E-18 puc = 5.994178352937092E-25 ud = 0
+ up = 0 lp = 1 eu = 1.67
+ vsat = 3.175301189774053E5 lvsat = -0.048910885952424 wvsat = -1.289675810099376
+ pvsat = 2.788787510213546E-7 a0 = 0.801114070626046 la0 = -4.975552000624815E-8
+ wa0 = 1.553459716743644E-6 pa0 = -3.672118569545672E-13 ags = 2.296937986912553
+ lags = -2.177505380219681E-7 wags = 1.483700385212299E-5 pags = -3.085918757195357E-12
+ b0 = 0 b1 = 1.560790734647861E-23 lb1 = -4.338810947432896E-30
+ wb1 = -1.090273542364144E-28 pb1 = 3.030829614947236E-35 keta = -0.257871825644216
+ lketa = 6.213763765233085E-8 wketa = 1.33287608886817E-8 pketa = -9.613594368509537E-14
+ a1 = 0 a2 = 0.806834430701736 la2 = -1.899889721914189E-9
+ wa2 = 5.395578782304452E-7 pa2 = -1.49990615453525E-13 rdsw = 547.88
+ rdswmin = 0 rdw = 0 rdwmin = 0
+ rsw = 0 rswmin = 0 prwb = -0.32348
+ prwg = 0.1376 wr = 1 voff = -0.120647836650487
+ lvoff = -3.838823789905296E-8 wvoff = 3.744690421810312E-7 pvoff = -1.13365531860351E-13
+ voffl = 0 minv = 0 nfactor = 2.159279675485483
+ lnfactor = -4.75324913110901E-8 wnfactor = -3.307498448344419E-6 pnfactor = 9.506658127697417E-13
+ eta0 = -4.454935738111374 leta0 = 9.481701072373007E-7 weta0 = 2.762053233900224E-5
+ peta0 = -5.647418335008352E-12 etab = 0.124971191967595 letab = -3.86474083082358E-8
+ wetab = 1.750962641995205E-7 petab = -3.115767794025613E-14 dsub = 0.917448105477036
+ ldsub = -1.423686095150368E-7 wdsub = -7.258647359483733E-7 pdsub = 2.237266145786823E-13
+ cit = 1E-5 cdsc = 1.3E-4 cdscb = 7.8E-4
+ cdscd = 0 pclm = 1.987077637342496 lpclm = -2.81622907551503E-7
+ wpclm = -5.655862716452216E-6 ppclm = 1.18119033511035E-12 pdiblc1 = 1.690366910248538
+ lpdiblc1 = -3.149170462851251E-7 wpdiblc1 = -3.965776888364217E-6 ppdiblc1 = 8.398712494523595E-13
+ pdiblc2 = 0.062510237832766 lpdiblc2 = -1.215658831985766E-8 wpdiblc2 = -2.433536578938812E-7
+ ppdiblc2 = 5.077730181243138E-14 pdiblcb = -0.569956859604857 lpdiblcb = 1.02945087315495E-7
+ wpdiblcb = 3.457467786420263E-6 ppdiblcb = -7.191118099619776E-13 drout = -4.009339495823783
+ ldrout = 1.051324274205383E-6 wdrout = 2.129990601077772E-5 pdrout = -4.569112177977646E-12
+ pscbe1 = 8E8 pscbe2 = -3.881242203276356E-8 lpscbe2 = 9.901447472260909E-15
+ wpscbe2 = 3.2653436561042E-13 ppscbe2 = -6.732346338218335E-20 pvag = 0
+ delta = 0.01 fprout = 0 pdits = 0
+ pditsl = 0 pditsd = 0 lambda = 0
+ vtl = 0 lc = 5E-9 xn = 3
+ alpha0 = 2.83319975417827E-8 lalpha0 = -5.8719167047203E-15 walpha0 = 2.577255956443585E-14
+ palpha0 = -5.360383118687884E-21 alpha1 = -2.971257142857143E-10 lalpha1 = 8.259738306285714E-17
+ beta0 = 35.96521863071619 lbeta0 = -5.679097758915601E-6 wbeta0 = 2.700163867911603E-6
+ pbeta0 = -6.415383425741376E-13 aigbacc = 0.43 bigbacc = 0.054
+ cigbacc = 0.075 nigbacc = 1 aigbinv = 0.35
+ bigbinv = 0.03 cigbinv = 6E-3 eigbinv = 1.1
+ nigbinv = 3 aigc = 0.43 bigc = 0.054
+ cigc = 0.075 aigsd = 0.43 bigsd = 0.054
+ cigsd = 0.075 dlcig = 0 nigc = 1
+ poxedge = 1 pigcd = 1 ntox = 1
+ toxref = 4.23E-9 agidl = -3.496829594150376E-11 lagidl = 3.751956665218676E-17
+ wagidl = 6.728698898340645E-16 pagidl = -1.87049754935192E-22 bgidl = 1.918143089397852E9
+ lbgidl = -239.2535925388794 wbgidl = 9.18719470873238E3 pbgidl = -1.573495742495903E-3
+ cgidl = -362.58942597944235 lcgidl = 1.378106495306122E-4 wcgidl = -1.863281528716099E-3
+ pcgidl = 3.875401985946041E-10 egidl = 0.1 noia = 1.5E42
+ noib = 0 noic = 0 em = 4.1E7
+ af = 1 ef = 1 kf = 0
+ lintnoi = -2E-7 tnoia = 2.5E7 tnoib = 0
+ ntnoi = 1 rnoia = 0.69 rnoib = 0.34
+ xpart = 0 cgso = {5.248925E-11/sw_func_tox_lv_ratio} cgdo = {5.248925E-11/sw_func_tox_lv_ratio}
+ cgbo = {0/sw_func_tox_lv_ratio} ckappas = 0.6 cf = 1.2E-11
+ clc = 1E-7 cle = 0.6 dlc = -3E-9
+ dwc = 0 vfbcv = -0.14469 noff = 3.9
+ voffcv = -0.10701 acde = 0.8 moin = 18.13
+ cgsl = {9.548271750000001E-12/sw_func_tox_lv_ratio} cgdl = {9.548271750000001E-12/sw_func_tox_lv_ratio} ijthsrev = 0.1
+ ijthsfwd = 0.1 xjbvs = 1 bvs = 12.69
+ jss = 2.1483E-5 jsws = 8.040000000000001E-10 cjs = {sw_psd_nw_cj}
+ mjs = 0.34629 mjsws = 0.29781 cjsws = {9.888891999999999E-11*sw_func_psd_nw_cj}
+ cjswgs = {2.39155046E-10*sw_func_psd_nw_cj} mjswgs = 0.9274 pbs = 0.6587
+ pbsws = 0.7418 pbswgs = 1.4338 xrcrg1 = 12
+ xrcrg2 = 1 rbpb = 50 rbpd = 50
+ rbps = 50 rbdb = 50 rbsb = 50
+ gbmin = 1E-12 tnom = 30 ute = -1.17383484310212
+ lute = 1.817471613471237E-7 wute = 4.356409410889532E-6 pute = -9.060808805520919E-13
+ kt1 = -0.53621646549 wkt1 = -1.584533850345847E-7 kt1l = 0
+ kt2 = -0.131083267726 wkt2 = 6.372960321171207E-8 ua1 = -1.985849578859898E-10
+ lua1 = 6.930263278079127E-17 wua1 = 2.327567313818122E-15 pua1 = -4.841060704664037E-22
+ ub1 = 2.371845547121538E-19 lub1 = 3.234534643452857E-26 wub1 = 1.086336378493248E-24
+ pub1 = -2.259449306900537E-31 uc1 = 9.504779912119998E-11 wuc1 = -3.986060318913972E-16
+ at = 6.127424664301832E5 lat = -0.12744072746493 wat = -2.655502897184643
+ pat = 6.075056570558788E-7 prt = 0 njs = 1.3632
+ xtis = 5.2 tpb = 2.0386E-3 tpbsw = 1.246E-3
+ tpbswg = 0 tcj = 1.2407E-3 tcjsw = 3.7357E-4
+ tcjswg = 2E-12 tvoff = 0 tvfbsdoff = 0
+ saref = 1.25E-6 sbref = 1.24E-6 wlod = 0
+ ku0 = 4.5E-8 kvsat = 0.5 kvth0 = 3.29E-8
+ tku0 = 0 llodku0 = 0 wlodku0 = 1
+ llodvth = 0 wlodvth = 1 lku0 = 0
+ wku0 = 2.5E-7 pku0 = 0 lkvth0 = 0
+ wkvth0 = 2E-7 pkvth0 = 0 stk2 = 0
+ lodk2 = 1 steta0 = 0 lodeta0 = 1

.model pshort_model.16 pmos
+ level = 54 lmin = 1.5E-7 lmax = 1.8E-7 wmin = 5E-6
+ wmax = 7E-6 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 4.23E-9
+ toxm = 4.23E-9 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 9.999999999999999E22 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {7.3039E-9+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {-1.3994E-8-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = -5.722E-9 dwb = -1.7864E-8 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = -0.851929258852923 lvth0 = -3.82222701405814E-8
+ wvth0 = -4.60082068110547E-8 pvth0 = 2.554757782774253E-14 k1 = -0.724663606244711
+ lk1 = 3.566574150976426E-7 wk1 = 1.171721054647535E-6 pk1 = -1.971267435011108E-13
+ k2 = 0.545043873773805 lk2 = -1.498589836171933E-7 wk2 = -4.512898020382907E-7
+ pk2 = 8.274493037395078E-14 k3 = -15.845 k3b = 2
+ w0 = 0 lpe0 = 0 lpeb = 0
+ vbm = -3 dvtp0 = 0 dvtp1 = 0
+ dvt0 = 4.4955 dvt1 = 0.294 dvt2 = 0.015
+ dvt0w = -4.9772 dvt1w = 1.1472E6 dvt2w = -8.96E-3
+ vfbsdoff = 0 u0 = 8.030755119963514E-3 lu0 = -8.110879611687108E-10
+ wu0 = -7.662534576663606E-9 pu0 = 1.015457130478545E-15 ua = -1.135672078347297E-9
+ lua = -2.393042182320217E-16 wua = 1.865991680551048E-15 pua = -3.694386025335525E-22
+ ub = 1.448674775370495E-18 lub = 1.404412514608591E-25 wub = -5.180478926431614E-24
+ pub = 9.922945662243082E-31 uc = -6.916243117904054E-13 luc = 1.427577615844065E-19
+ wuc = 6.909949140157484E-18 puc = -1.204247714375102E-24 ud = 0
+ up = 0 lp = 1 eu = 1.67
+ vsat = 3.373885035051632E5 lvsat = -0.053041191633583 wvsat = -0.42236335745069
+ pvsat = 9.848816861985972E-8 a0 = 1.287211766853238 la0 = -1.508580076491492E-7
+ wa0 = -1.675177245749992E-5 pa0 = 3.440056772502004E-12 ags = 1.25
+ b0 = 0 b1 = -3.641845047511675E-23 lb1 = 6.482047163165079E-30
+ wb1 = 2.543971598849668E-28 pb1 = -4.527964169360547E-35 keta = 0.326538314613292
+ lketa = -5.941265859954758E-8 wketa = -3.035757967665067E-6 pketa = 5.380375068133416E-13
+ a1 = 0 a2 = -2.889952837126629 la2 = 7.669875005391718E-7
+ wa2 = 1.613735198731628E-5 pa2 = -3.394144616614069E-12 rdsw = 547.88
+ rdswmin = 0 rdw = 0 rdwmin = 0
+ rsw = 0 rswmin = 0 prwb = -0.32348
+ prwg = 0.1376 wr = 1 voff = 0.158821789465681
+ lvoff = -9.651456649570254E-8 wvoff = -8.575431171881143E-7 pvoff = 1.428782131425188E-13
+ voffl = 0 minv = 0 nfactor = -0.950436192991012
+ lnfactor = 5.992510927415992E-7 wnfactor = 6.495771677716697E-6 pnfactor = -1.088296734209458E-12
+ eta0 = -1.897520054157942 leta0 = 4.162583339631943E-7 weta0 = 7.612484234703244E-6
+ peta0 = -1.485984425891413E-12 etab = -0.272547274226358 letab = 4.403166243851222E-8
+ wetab = -1.41635294846011E-7 petab = 3.471868556250587E-14 dsub = 0.072423568230697
+ ldsub = 3.338635393775472E-8 wdsub = 2.425181995941734E-6 pdsub = -4.316532930936773E-13
+ cit = 1E-5 cdsc = 1.3E-4 cdscb = 7.8E-4
+ cdscd = 0 pclm = 4.439190831633557 lpclm = -7.916330266057121E-7
+ wpclm = -1.371199229420316E-5 ppclm = 2.856768613727612E-12 pdiblc1 = 1.10627484963891
+ lpdiblc1 = -1.9343290678305E-7 wpdiblc1 = 5.012357479854526E-7 ppdiblc1 = -8.921377475673567E-14
+ pdiblc2 = 0.041029720268646 lpdiblc2 = -7.68889843273149E-9 wpdiblc2 = -1.023009550259961E-7
+ ppdiblc2 = 2.144003224834569E-14 pdiblcb = -1.565240203789704 lpdiblcb = 3.099520795058129E-7
+ wpdiblcb = 7.429431888099599E-6 ppdiblcb = -1.545232679542059E-12 drout = 1.314725704932861
+ ldrout = -5.601739876959001E-8 wdrout = -4.632910886933662E-6 pdrout = 8.246025429435486E-13
+ pscbe1 = 1.091897231410302E9 lpscbe1 = -60.71112136656592 wpscbe1 = -1.455222180674515E3
+ ppscbe1 = 3.02668750914131E-4 pscbe2 = 1.20890865910322E-8 lpscbe2 = -6.854555033851235E-16
+ wpscbe2 = -1.208873650157495E-14 ppscbe2 = 3.10607837988625E-21 pvag = 0
+ delta = 0.01 fprout = 0 pdits = 0
+ pditsl = 0 pditsd = 0 lambda = 0
+ vtl = 0 lc = 5E-9 xn = 3
+ alpha0 = 1E-10 alpha1 = 1E-10 beta0 = 21.02500547532119
+ lbeta0 = -2.571712705151307E-6 wbeta0 = -3.585736170584074E-5 pbeta0 = 7.377964286459464E-12
+ aigbacc = 0.43 bigbacc = 0.054 cigbacc = 0.075
+ nigbacc = 1 aigbinv = 0.35 bigbinv = 0.03
+ cigbinv = 6E-3 eigbinv = 1.1 nigbinv = 3
+ aigc = 0.43 bigc = 0.054 cigc = 0.075
+ aigsd = 0.43 bigsd = 0.054 cigsd = 0.075
+ dlcig = 0 nigc = 1 poxedge = 1
+ pigcd = 1 ntox = 1 toxref = 4.23E-9
+ agidl = 9.947975291485523E-10 lagidl = -1.766593677766438E-16 wagidl = -5.620659632966552E-15
+ pagidl = 1.121928863453063E-21 bgidl = -1.559685729112315E9 lbgidl = 484.0930677654131
+ wbgidl = 1.598042711244777E4 pbgidl = -2.98640656367986E-3 cgidl = 300
+ egidl = 0.1 noia = 1.5E42 noib = 0
+ noic = 0 em = 4.1E7 af = 1
+ ef = 1 kf = 0 lintnoi = -2E-7
+ tnoia = 2.5E7 tnoib = 0 ntnoi = 1
+ rnoia = 0.69 rnoib = 0.34 xpart = 0
+ cgso = {5.248925E-11/sw_func_tox_lv_ratio} cgdo = {5.248925E-11/sw_func_tox_lv_ratio} cgbo = {0/sw_func_tox_lv_ratio}
+ ckappas = 0.6 cf = 1.2E-11 clc = 1E-7
+ cle = 0.6 dlc = -3E-9 dwc = 0
+ vfbcv = -0.14469 noff = 3.9 voffcv = -0.10701
+ acde = 0.8 moin = 18.13 cgsl = {9.548271750000001E-12/sw_func_tox_lv_ratio}
+ cgdl = {9.548271750000001E-12/sw_func_tox_lv_ratio} ijthsrev = 0.1 ijthsfwd = 0.1
+ xjbvs = 1 bvs = 12.69 jss = 2.1483E-5
+ jsws = 8.040000000000001E-10 cjs = {sw_psd_nw_cj} mjs = 0.34629
+ mjsws = 0.29781 cjsws = {9.888891999999999E-11*sw_func_psd_nw_cj} cjswgs = {2.39155046E-10*sw_func_psd_nw_cj}
+ mjswgs = 0.9274 pbs = 0.6587 pbsws = 0.7418
+ pbswgs = 1.4338 xrcrg1 = 12 xrcrg2 = 1
+ rbpb = 50 rbpd = 50 rbps = 50
+ rbdb = 50 rbsb = 50 gbmin = 1E-12
+ tnom = 30 ute = -0.3 kt1 = 0.331803993177515
+ lkt1 = -1.805378391573392E-7 wkt1 = -7.886258637260403E-7 pkt1 = 1.310683134980785E-13
+ kt1l = 0 kt2 = -0.18521100692651 lkt2 = 1.125792022083557E-8
+ wkt2 = 4.418330904265854E-7 pkt2 = -7.864098809884708E-14 ua1 = 1.3462E-10
+ ub1 = 3.927E-19 uc1 = 4.335975821206713E-10 luc1 = -7.041429226649401E-17
+ wuc1 = -2.763509045367596E-15 puc1 = 4.918714479668877E-22 at = -2.253730452349742E5
+ lat = 0.046877241575283 wat = 1.839764015874636 pat = -3.274559176574947E-7
+ prt = 0 njs = 1.3632 xtis = 5.2
+ tpb = 2.0386E-3 tpbsw = 1.246E-3 tpbswg = 0
+ tcj = 1.2407E-3 tcjsw = 3.7357E-4 tcjswg = 2E-12
+ tvoff = 0 tvfbsdoff = 0 saref = 1.1E-6
+ sbref = 1.1E-6 wlod = 0 ku0 = 4.5E-8
+ kvsat = 0.5 kvth0 = 3.29E-8 tku0 = 0
+ llodku0 = 0 wlodku0 = 1 llodvth = 0
+ wlodvth = 1 lku0 = 0 wku0 = 2.5E-7
+ pku0 = 0 lkvth0 = 0 wkvth0 = 2E-7
+ pkvth0 = 0 stk2 = 0 lodk2 = 1
+ steta0 = 0 lodeta0 = 1

.model pshort_model.17 pmos
+ level = 54 lmin = 8E-6 lmax = 2.02E-5 wmin = 3E-6
+ wmax = 5E-6 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 4.23E-9
+ toxm = 4.23E-9 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 9.999999999999999E22 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {7.3039E-9+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {-1.3994E-8-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = -5.722E-9 dwb = -1.7864E-8 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = -1.065871703871769 wvth0 = 5.402128049618837E-8
+ k1 = 0.44180966168701 wk1 = -5.606632733867083E-8 k2 = 0.021576800612952
+ wk2 = -6.631649116398325E-10 k3 = -15.845 k3b = 2
+ w0 = 0 lpe0 = 0 lpeb = 0
+ vbm = -3 dvtp0 = 0 dvtp1 = 0
+ dvt0 = 4.4955 dvt1 = 0.294 dvt2 = 0.015
+ dvt0w = -4.9772 dvt1w = 1.1472E6 dvt2w = -8.96E-3
+ vfbsdoff = 0 u0 = 8.560047547549998E-3 wu0 = 8.963498132415108E-9
+ ua = -1.096266560575684E-9 wua = 2.69429165360946E-15 ub = 1.234728874152449E-18
+ wub = -1.52418976106254E-24 uc = -1.04160361652318E-11 wuc = -2.632876845259807E-16
+ ud = 0 up = 0 lp = 1
+ eu = 1.67 vsat = 3.1984364933945E5 wvsat = -0.795325347573929
+ a0 = 1.3212940808532 wa0 = -6.326317170883117E-7 ags = 0.296239212736026
+ wags = -3.408782991798867E-7 b0 = 0 b1 = 0
+ keta = -0.012125816957524 wketa = 3.621515900697344E-8 a1 = 0
+ a2 = 1.073632922557868 wa2 = -8.169015926674631E-7 rdsw = 547.88
+ rdswmin = 0 rdw = 0 rdwmin = 0
+ rsw = 0 rswmin = 0 prwb = -0.32348
+ prwg = 0.1376 wr = 1 voff = -0.251471733730319
+ wvoff = -3.238691591704484E-9 voffl = 0 minv = 0
+ nfactor = 1.28816711935094 wnfactor = 1.363870099476235E-6 eta0 = 0.08
+ etab = -0.07 dsub = 0.56 cit = 1E-5
+ cdsc = 1.3E-4 cdscb = 7.8E-4 cdscd = 0
+ pclm = 0.344479425579197 wpclm = -5.842665564680252E-7 pdiblc1 = 0.39
+ pdiblc2 = 1.34084551929727E-4 wpdiblc2 = 1.725719337864981E-10 pdiblcb = -0.025
+ drout = 0.56 pscbe1 = 8.63994449244292E8 wpscbe1 = -319.0374281057893
+ pscbe2 = 7.8886136971903E-9 wpscbe2 = 5.924890869715114E-15 pvag = 0
+ delta = 0.01 fprout = 0 pdits = 0
+ pditsl = 0 pditsd = 0 lambda = 0
+ vtl = 0 lc = 5E-9 xn = 3
+ alpha0 = 2.226759885480409E-10 walpha0 = -6.115879164346925E-16 alpha1 = 2.492695158757741E-10
+ walpha1 = -7.441670801448602E-16 beta0 = 1.382664626227562 wbeta0 = 2.476991752517078E-5
+ aigbacc = 0.43 bigbacc = 0.054 cigbacc = 0.075
+ nigbacc = 1 aigbinv = 0.35 bigbinv = 0.03
+ cigbinv = 6E-3 eigbinv = 1.1 nigbinv = 3
+ aigc = 0.43 bigc = 0.054 cigc = 0.075
+ aigsd = 0.43 bigsd = 0.054 cigsd = 0.075
+ dlcig = 0 nigc = 1 poxedge = 1
+ pigcd = 1 ntox = 1 toxref = 4.23E-9
+ agidl = 1E-10 bgidl = 1.82580602497249E9 wbgidl = -1.412883206781777E3
+ cgidl = 300 egidl = 0.1 noia = 1.5E42
+ noib = 0 noic = 0 em = 4.1E7
+ af = 1 ef = 1 kf = 0
+ lintnoi = -2E-7 tnoia = 2.5E7 tnoib = 0
+ ntnoi = 1 rnoia = 0.69 rnoib = 0.34
+ xpart = 0 cgso = {5.248925E-11/sw_func_tox_lv_ratio} cgdo = {5.248925E-11/sw_func_tox_lv_ratio}
+ cgbo = {0/sw_func_tox_lv_ratio} ckappas = 0.6 cf = 1.2E-11
+ clc = 1E-7 cle = 0.6 dlc = -3E-9
+ dwc = 0 vfbcv = -0.14469 noff = 3.9
+ voffcv = -0.10701 acde = 0.8 moin = 18.13
+ cgsl = {9.548271750000001E-12/sw_func_tox_lv_ratio} cgdl = {9.548271750000001E-12/sw_func_tox_lv_ratio} ijthsrev = 0.1
+ ijthsfwd = 0.1 xjbvs = 1 bvs = 12.69
+ jss = 2.1483E-5 jsws = 8.040000000000001E-10 cjs = {sw_psd_nw_cj}
+ mjs = 0.34629 mjsws = 0.29781 cjsws = {9.888891999999999E-11*sw_func_psd_nw_cj}
+ cjswgs = {2.39155046E-10*sw_func_psd_nw_cj} mjswgs = 0.9274 pbs = 0.6587
+ pbsws = 0.7418 pbswgs = 1.4338 xrcrg1 = 12
+ xrcrg2 = 1 rbpb = 50 rbpd = 50
+ rbps = 50 rbdb = 50 rbsb = 50
+ gbmin = 1E-12 tnom = 30 ute = -0.154965580668972
+ wute = -4.859027130397824E-8 kt1 = -0.423714028857974 wkt1 = -6.151780113848939E-8
+ kt1l = 0 kt2 = -0.047357787652513 wkt2 = -1.58429699261116E-8
+ ua1 = 1.73469673296457E-9 wua1 = 1.120019044389131E-15 ub1 = -7.732550472225199E-19
+ wub1 = 1.038351865016307E-25 uc1 = 1.1392027463169E-10 wuc1 = -9.919009265833227E-18
+ at = 9E4 prt = 0 njs = 1.3632
+ xtis = 5.2 tpb = 2.0386E-3 tpbsw = 1.246E-3
+ tpbswg = 0 tcj = 1.2407E-3 tcjsw = 3.7357E-4
+ tcjswg = 2E-12 tvoff = 0 tvfbsdoff = 0
+ saref = 3E-6 sbref = 3E-6 wlod = 0
+ ku0 = 4.5E-8 kvsat = 0.5 kvth0 = 3.29E-8
+ tku0 = 0 llodku0 = 0 wlodku0 = 1
+ llodvth = 0 wlodvth = 1 lku0 = 0
+ wku0 = 2.5E-7 pku0 = 0 lkvth0 = 0
+ wkvth0 = 2E-7 pkvth0 = 0 stk2 = 0
+ lodk2 = 1 steta0 = 0 lodeta0 = 1

.model pshort_model.18 pmos
+ level = 54 lmin = 4E-6 lmax = 8E-6 wmin = 3E-6
+ wmax = 5E-6 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 4.23E-9
+ toxm = 4.23E-9 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 9.999999999999999E22 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {7.3039E-9+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {-1.3994E-8-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = -5.722E-9 dwb = -1.7864E-8 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = -1.069634370512243 lvth0 = 3.020664263772474E-8
+ wvth0 = 5.046909553994925E-8 pvth0 = 2.85168982024682E-14 k1 = 0.52976404061942
+ lk1 = -7.060966986168385E-7 wk1 = -4.16088763066334E-7 pk1 = 2.890255793752451E-12
+ k2 = -0.010211893465789 lk2 = 2.551992545998025E-7 wk2 = 1.324597585732309E-7
+ pk2 = -1.06870923226146E-12 k3 = -15.845 k3b = 2
+ w0 = 0 lpe0 = 0 lpeb = 0
+ vbm = -3 dvtp0 = 0 dvtp1 = 0
+ dvt0 = 4.4955 dvt1 = 0.294 dvt2 = 0.015
+ dvt0w = -4.9772 dvt1w = 1.1472E6 dvt2w = -8.96E-3
+ vfbsdoff = 0 u0 = 6.294102812122239E-3 lu0 = 1.819097714467722E-8
+ wu0 = 1.650445362260968E-8 pu0 = -6.053870018381617E-14 ua = -1.630667962144931E-9
+ lua = 4.290168038981094E-15 wua = 4.56788547139998E-15 pua = -1.504118868609647E-20
+ ub = 1.545456020208192E-18 lub = -2.494513799809752E-24 wub = -2.613424091440998E-24
+ pub = 8.744360133466297E-30 uc = 4.582367216757989E-12 luc = -1.204070023697733E-16
+ wuc = -3.482631921330051E-16 puc = 6.821823553631002E-22 ud = 0
+ up = 0 lp = 1 eu = 1.67
+ vsat = 5.442673188696277E5 lvsat = -1.801670525904231 wvsat = -1.394322094091133
+ pvsat = 4.808738693079152E-6 a0 = 1.338105178974543 la0 = -1.349592939849679E-7
+ wa0 = -6.328490356903333E-7 pa0 = 1.744631129206658E-15 ags = 0.334396635782315
+ lags = -3.063273343265348E-7 wags = -9.525074912703755E-7 pags = 4.910151814552139E-12
+ b0 = 0 b1 = 0 keta = -0.012690290320559
+ lketa = 4.53158538476452E-9 wketa = 6.704534538456111E-8 pketa = -2.475043662770373E-13
+ a1 = 0 a2 = 1.349180454674873 la2 = -2.212092281264934E-6
+ wa2 = -1.639519045778821E-6 pa2 = 6.603963042168541E-12 rdsw = 547.88
+ rdswmin = 0 rdw = 0 rdwmin = 0
+ rsw = 0 rswmin = 0 prwb = -0.32348
+ prwg = 0.1376 wr = 1 voff = -0.253832649645215
+ lvoff = 1.895340463379359E-8 wvoff = 9.254325728505738E-10 pvoff = -3.342953882355803E-14
+ voffl = 0 minv = 0 nfactor = 1.223183052665572
+ lnfactor = 5.21691307541335E-7 wnfactor = 1.727037959687108E-6 pnfactor = -2.915507223758564E-12
+ eta0 = 0.08 etab = -0.07 dsub = 0.56
+ cit = 1E-5 cdsc = 1.3E-4 cdscb = 7.8E-4
+ cdscd = 0 pclm = 0.206725750144198 lpclm = 1.105884853348064E-6
+ wpclm = -9.665104936895698E-7 ppclm = 3.068649741087312E-12 pdiblc1 = 0.39
+ pdiblc2 = 3.22442719140064E-4 lpdiblc2 = -1.512137106066579E-9 wpdiblc2 = -4.592262230704906E-10
+ ppdiblc2 = 5.072068021670023E-15 pdiblcb = -0.025 drout = 0.56
+ pscbe1 = 9.284366676499462E8 lpscbe1 = -517.3413560539722 wpscbe1 = -640.3071610960347
+ ppscbe1 = 2.579149561208895E-3 pscbe2 = 6.369823655948436E-9 lpscbe2 = 1.219282822560919E-14
+ wpscbe2 = 1.154737197936684E-14 ppscbe2 = -4.513721087851072E-20 pvag = 0
+ delta = 0.01 fprout = 0 pdits = 0
+ pditsl = 0 pditsd = 0 lambda = 0
+ vtl = 0 lc = 5E-9 xn = 3
+ alpha0 = 2.1778265896932E-10 lalpha0 = 3.928359113801638E-17 walpha0 = -5.87192749320908E-16
+ palpha0 = -1.958441088474562E-22 alpha1 = 2.506003080151116E-10 lalpha1 = -1.068358332509598E-17
+ walpha1 = -7.508016008961347E-16 palpha1 = 5.326185297698333E-23 beta0 = -9.458283719412403
+ lbeta0 = 8.703100322741752E-5 wbeta0 = 7.721546820757105E-5 pbeta0 = -4.210322515317011E-10
+ aigbacc = 0.43 bigbacc = 0.054 cigbacc = 0.075
+ nigbacc = 1 aigbinv = 0.35 bigbinv = 0.03
+ cigbinv = 6E-3 eigbinv = 1.1 nigbinv = 3
+ aigc = 0.43 bigc = 0.054 cigc = 0.075
+ aigsd = 0.43 bigsd = 0.054 cigsd = 0.075
+ dlcig = 0 nigc = 1 poxedge = 1
+ pigcd = 1 ntox = 1 toxref = 4.23E-9
+ agidl = 1.537202721633743E-10 lagidl = -4.312657002843023E-16 wagidl = -2.67816625825163E-16
+ pagidl = 2.150028658324898E-21 bgidl = 1.435872467176342E9 lbgidl = 3.130381922784789E3
+ wbgidl = 811.0571982624068 pbgidl = -0.01785376688441 cgidl = 300
+ egidl = 0.1 noia = 1.5E42 noib = 0
+ noic = 0 em = 4.1E7 af = 1
+ ef = 1 kf = 0 lintnoi = -2E-7
+ tnoia = 2.5E7 tnoib = 0 ntnoi = 1
+ rnoia = 0.69 rnoib = 0.34 xpart = 0
+ cgso = {5.248925E-11/sw_func_tox_lv_ratio} cgdo = {5.248925E-11/sw_func_tox_lv_ratio} cgbo = {0/sw_func_tox_lv_ratio}
+ ckappas = 0.6 cf = 1.2E-11 clc = 1E-7
+ cle = 0.6 dlc = -3E-9 dwc = 0
+ vfbcv = -0.14469 noff = 3.9 voffcv = -0.10701
+ acde = 0.8 moin = 18.13 cgsl = {9.548271750000001E-12/sw_func_tox_lv_ratio}
+ cgdl = {9.548271750000001E-12/sw_func_tox_lv_ratio} ijthsrev = 0.1 ijthsfwd = 0.1
+ xjbvs = 1 bvs = 12.69 jss = 2.1483E-5
+ jsws = 8.040000000000001E-10 cjs = {sw_psd_nw_cj} mjs = 0.34629
+ mjsws = 0.29781 cjsws = {9.888891999999999E-11*sw_func_psd_nw_cj} cjswgs = {2.39155046E-10*sw_func_psd_nw_cj}
+ mjswgs = 0.9274 pbs = 0.6587 pbsws = 0.7418
+ pbswgs = 1.4338 xrcrg1 = 12 xrcrg2 = 1
+ rbpb = 50 rbpd = 50 rbps = 50
+ rbdb = 50 rbsb = 50 gbmin = 1E-12
+ tnom = 30 ute = -0.02882875949875 lute = -1.01262488671269E-6
+ wute = -4.72207773603336E-7 pute = 3.400796225049216E-12 kt1 = -0.36925500460282
+ lkt1 = -4.371963932120831E-7 wkt1 = -1.98403491304958E-7 pkt1 = 1.098916678028128E-12
+ kt1l = 0 kt2 = -0.043259497821033 lkt2 = -3.290102158764008E-8
+ wkt2 = -3.179679311279622E-8 pkt2 = 1.280771010968258E-13 ua1 = 1.284925684797492E-9
+ lua1 = 3.610756577432718E-15 wua1 = 2.247874862031854E-15 pua1 = -9.054412969765964E-21
+ ub1 = -6.222704356621359E-19 lub1 = -1.212102649791425E-24 wub1 = 2.083969078032133E-25
+ pub1 = -8.394202438684493E-31 uc1 = 3.59891340229908E-10 luc1 = -1.974652762969706E-15
+ wuc1 = -1.99074218394995E-17 puc1 = 8.018685628044188E-23 at = 1.349728711382837E4
+ lat = 0.614162861017631 wat = 0.359699755072383 pat = -2.88766531732403E-6
+ prt = 0 njs = 1.3632 xtis = 5.2
+ tpb = 2.0386E-3 tpbsw = 1.246E-3 tpbswg = 0
+ tcj = 1.2407E-3 tcjsw = 3.7357E-4 tcjswg = 2E-12
+ tvoff = 0 tvfbsdoff = 0 saref = 3E-6
+ sbref = 3E-6 wlod = 0 ku0 = 4.5E-8
+ kvsat = 0.5 kvth0 = 3.29E-8 tku0 = 0
+ llodku0 = 0 wlodku0 = 1 llodvth = 0
+ wlodvth = 1 lku0 = 0 wku0 = 2.5E-7
+ pku0 = 0 lkvth0 = 0 wkvth0 = 2E-7
+ pkvth0 = 0 stk2 = 0 lodk2 = 1
+ steta0 = 0 lodeta0 = 1

.model pshort_model.19 pmos
+ level = 54 lmin = 2E-6 lmax = 4E-6 wmin = 3E-6
+ wmax = 5E-6 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 4.23E-9
+ toxm = 4.23E-9 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 9.999999999999999E22 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {7.3039E-9+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {-1.3994E-8-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = -5.722E-9 dwb = -1.7864E-8 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = -1.07232599320665 lvth0 = 4.104846655132381E-8
+ wvth0 = 6.503430675832252E-8 pvth0 = -3.015159780260476E-14 k1 = 0.37366012860566
+ lk1 = -7.731201427235578E-8 wk1 = 6.930740703625549E-8 pk1 = 9.350858453332617E-13
+ k2 = 0.044901793324714 lk2 = 3.320198557189578E-8 wk2 = -4.367877804313092E-8
+ pk2 = -3.592253204331943E-13 k3 = -15.845 k3b = 2
+ w0 = 0 lpe0 = 0 lpeb = 0
+ vbm = -3 dvtp0 = 0 dvtp1 = 0
+ dvt0 = 4.4955 dvt1 = 0.294 dvt2 = 0.015
+ dvt0w = -4.9772 dvt1w = 1.1472E6 dvt2w = -8.96E-3
+ vfbsdoff = 0 u0 = 0.01365820131878 lu0 = -1.147152327095725E-8
+ wu0 = -2.365863724033549E-11 pu0 = 6.036337661512589E-15 ua = 1.350736312895203E-10
+ lua = -2.822217910473754E-15 wua = 3.063364528058157E-16 pua = 2.124279622212597E-21
+ ub = 4.632524910383536E-19 lub = 1.864589029244009E-24 wub = 1.172412585385551E-25
+ pub = -2.254727128267146E-30 uc = -6.163134734900565E-11 luc = 1.463010453365479E-16
+ wuc = -1.332157545928835E-16 puc = -1.840261424792589E-22 ud = 0
+ up = 0 lp = 1 eu = 1.67
+ vsat = 9.750357883221177E4 lvsat = -2.111542198400747E-3 wvsat = -0.186289436856035
+ pvsat = -5.720235387193636E-8 a0 = 1.117324081705906 la0 = 7.543443164399372E-7
+ wa0 = 4.191536808280222E-7 pa0 = -4.235709686974131E-12 ags = 0.255210029904591
+ lags = 1.263536390966903E-8 wags = -4.71617893853999E-7 pags = 2.973134286834143E-12
+ b0 = 0 b1 = 0 keta = -0.013943011735425
+ lketa = 9.57753221118938E-9 wketa = 4.931706144605436E-8 pketa = -1.760950513121394E-13
+ a1 = 0 a2 = 0.8 rdsw = 547.88
+ rdswmin = 0 rdw = 0 rdwmin = 0
+ rsw = 0 rswmin = 0 prwb = -0.32348
+ prwg = 0.1376 wr = 1 voff = -0.245204931884238
+ lvoff = -1.579893897480877E-8 wvoff = -4.33580592351116E-8 pvoff = 1.449438347770119E-13
+ voffl = 0 minv = 0 nfactor = 1.674555738855786
+ lnfactor = -1.296432455960615E-6 wnfactor = 3.733757940830673E-7 pnfactor = 2.537027735348525E-12
+ eta0 = 0.280942516865585 leta0 = -8.093940466243725E-7 weta0 = -5.998922224988847E-7
+ peta0 = 2.416358673518838E-12 etab = -0.245666731739443 letab = 7.075834874456966E-7
+ wetab = 5.244340907344263E-7 petab = -2.112414224269181E-12 dsub = 1.31827366676702
+ ldsub = -3.054317230453556E-6 wdsub = -2.263744290231661E-6 pdsub = 9.11833483612165E-12
+ cit = 1E-5 cdsc = 1.3E-4 cdscb = 7.8E-4
+ cdscd = 0 pclm = -0.016710752485446 lpclm = 2.005884404702241E-6
+ wpclm = 1.272727704465195E-6 ppclm = -5.950974850221704E-12 pdiblc1 = 0.39
+ pdiblc2 = -8.681090225245465E-4 lpdiblc2 = 3.283391022737572E-9 wpdiblc2 = 3.233505227594406E-9
+ ppdiblc2 = -9.80220994883077E-15 pdiblcb = 0.010814953456534 lpdiblcb = -1.442622027434792E-7
+ wpdiblcb = -1.785515896055698E-7 ppdiblcb = 7.192036603121599E-13 drout = 0.56
+ pscbe1 = 8.291911349705855E8 lpscbe1 = -117.5815413678988 wpscbe1 = -87.14698665033322
+ ppscbe1 = 3.510270164637024E-4 pscbe2 = 8.699702033138665E-9 lpscbe2 = 2.808106080827472E-15
+ wpscbe2 = 3.869622743212853E-15 ppscbe2 = -1.42113290882733E-20 pvag = 0
+ delta = 0.01 fprout = 0 pdits = 0
+ pditsl = 0 pditsd = 0 lambda = 0
+ vtl = 0 lc = 5E-9 xn = 3
+ alpha0 = 2.818313550153944E-10 lalpha0 = -2.187037879512186E-16 walpha0 = -9.06500619009178E-16
+ palpha0 = 1.090324158562459E-21 alpha1 = 3.979663250780386E-10 lalpha1 = -6.042721316623615E-16
+ walpha1 = -1.485478992906718E-15 palpha1 = 3.01253357186691E-21 beta0 = 13.5215377181067
+ lbeta0 = -5.531441765052186E-6 wbeta0 = -4.205677710282384E-5 pbeta0 = 5.939492131162576E-11
+ aigbacc = 0.43 bigbacc = 0.054 cigbacc = 0.075
+ nigbacc = 1 aigbinv = 0.35 bigbinv = 0.03
+ cigbinv = 6E-3 eigbinv = 1.1 nigbinv = 3
+ aigc = 0.43 bigc = 0.054 cigc = 0.075
+ aigsd = 0.43 bigsd = 0.054 cigsd = 0.075
+ dlcig = 0 nigc = 1 poxedge = 1
+ pigcd = 1 ntox = 1 toxref = 4.23E-9
+ agidl = 8.17290400784875E-11 lagidl = -1.412858813411635E-16 wagidl = 9.108790107922108E-17
+ pagidl = 7.04365530808362E-22 bgidl = 2.570451567502817E9 lbgidl = -1.439689078381049E3
+ wbgidl = -4.688413860100682E3 pbgidl = 4.298036545023972E-3 cgidl = 300
+ egidl = 0.1 noia = 1.5E42 noib = 0
+ noic = 0 em = 4.1E7 af = 1
+ ef = 1 kf = 0 lintnoi = -2E-7
+ tnoia = 2.5E7 tnoib = 0 ntnoi = 1
+ rnoia = 0.69 rnoib = 0.34 xpart = 0
+ cgso = {5.248925E-11/sw_func_tox_lv_ratio} cgdo = {5.248925E-11/sw_func_tox_lv_ratio} cgbo = {0/sw_func_tox_lv_ratio}
+ ckappas = 0.6 cf = 1.2E-11 clc = 1E-7
+ cle = 0.6 dlc = -3E-9 dwc = 0
+ vfbcv = -0.14469 noff = 3.9 voffcv = -0.10701
+ acde = 0.8 moin = 18.13 cgsl = {9.548271750000001E-12/sw_func_tox_lv_ratio}
+ cgdl = {9.548271750000001E-12/sw_func_tox_lv_ratio} ijthsrev = 0.1 ijthsfwd = 0.1
+ xjbvs = 1 bvs = 12.69 jss = 2.1483E-5
+ jsws = 8.040000000000001E-10 cjs = {sw_psd_nw_cj} mjs = 0.34629
+ mjsws = 0.29781 cjsws = {9.888891999999999E-11*sw_func_psd_nw_cj} cjswgs = {2.39155046E-10*sw_func_psd_nw_cj}
+ mjswgs = 0.9274 pbs = 0.6587 pbsws = 0.7418
+ pbswgs = 1.4338 xrcrg1 = 12 xrcrg2 = 1
+ rbpb = 50 rbpd = 50 rbps = 50
+ rbdb = 50 rbsb = 50 gbmin = 1E-12
+ tnom = 30 ute = -1.404237048321661 lute = 4.52750319576653E-6
+ wute = 6.42644637334934E-6 pute = -2.43868998950264E-11 kt1 = -0.50460799020204
+ lkt1 = 1.080038085457474E-7 wkt1 = 2.203432957900199E-7 pkt1 = -5.877903554289979E-13
+ kt1l = 0 kt2 = -0.075404117653803 lkt2 = 9.65771213633198E-8
+ wkt2 = 8.60291949947026E-8 pkt2 = -3.465245650883221E-13 ua1 = 3.369892806423134E-10
+ lua1 = 7.429033038132929E-15 wua1 = 1.264180075774855E-14 pua1 = -5.092102175060208E-20
+ ub1 = 4.581427676634733E-19 lub1 = -5.563994067828539E-24 wub1 = -8.779247296099418E-24
+ pub1 = 3.53627027577209E-29 uc1 = -5.355456819275394E-10 luc1 = 1.632156817036226E-15
+ wuc1 = 7.845429157980095E-16 puc1 = -3.160129450319393E-21 at = 1.744206800827801E5
+ lat = -0.034034634780591 wat = -0.324619589651941 pat = -1.312352086065888E-7
+ prt = 0 njs = 1.3632 xtis = 5.2
+ tpb = 2.0386E-3 tpbsw = 1.246E-3 tpbswg = 0
+ tcj = 1.2407E-3 tcjsw = 3.7357E-4 tcjswg = 2E-12
+ tvoff = 0 tvfbsdoff = 0 saref = 3E-6
+ sbref = 3E-6 wlod = 0 ku0 = 4.5E-8
+ kvsat = 0.5 kvth0 = 3.29E-8 tku0 = 0
+ llodku0 = 0 wlodku0 = 1 llodvth = 0
+ wlodvth = 1 lku0 = 0 wku0 = 2.5E-7
+ pku0 = 0 lkvth0 = 0 wkvth0 = 2E-7
+ pkvth0 = 0 stk2 = 0 lodk2 = 1
+ steta0 = 0 lodeta0 = 1

.model pshort_model.20 pmos
+ level = 54 lmin = 1E-6 lmax = 2E-6 wmin = 3E-6
+ wmax = 5E-6 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 4.23E-9
+ toxm = 4.23E-9 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 9.999999999999999E22 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {7.3039E-9+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {-1.3994E-8-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = -5.722E-9 dwb = -1.7864E-8 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = -1.054281269474241 lvth0 = 4.453983358684258E-9
+ wvth0 = -8.184980312001091E-9 pvth0 = 1.183362377445667E-13 k1 = 0.09806534196671
+ lk1 = 4.815909058939933E-7 wk1 = 1.338847399218746E-6 pk1 = -1.639526024332922E-12
+ k2 = 0.154627916744053 lk2 = -1.89321276009043E-7 wk2 = -5.433761550134114E-7
+ pk2 = 6.541549636940107E-13 k3 = -15.845 k3b = 2
+ w0 = 0 lpe0 = 0 lpeb = 0
+ vbm = -3 dvtp0 = 0 dvtp1 = 0
+ dvt0 = 4.4955 dvt1 = 0.294 dvt2 = 0.015
+ dvt0w = -4.9772 dvt1w = 1.1472E6 dvt2w = -8.96E-3
+ vfbsdoff = 0 u0 = 6.111550817111351E-3 lu0 = 3.832993386620291E-9
+ wu0 = 1.579483311776885E-8 pu0 = -2.604337379574497E-14 ua = -1.729783114022036E-9
+ lua = 9.596891907371398E-16 wua = 4.467019700126177E-15 pua = -6.313536075154129E-21
+ ub = 1.689397095498835E-18 lub = -6.220175148665935E-25 wub = -2.894828047246827E-24
+ pub = 3.85371327903394E-30 uc = 5.258435523131327E-11 luc = -8.532702890790793E-17
+ wuc = -4.551757686381062E-16 puc = 4.689049024842841E-22 ud = 0
+ up = 0 lp = 1 eu = 1.67
+ vsat = 2.44870871758392E5 lvsat = -0.300970643845179 wvsat = -0.823819744891491
+ pvsat = 1.235701460460272E-6 a0 = 2.853730841489874 la0 = -2.767067755520834E-6
+ wa0 = -6.115946966166749E-6 pa0 = 9.0173960039235E-12 ags = -1.466879113629511
+ lags = 3.505011481927105E-6 wags = 6.013220331301E-6 pags = -1.017803981572149E-11
+ b0 = 0 b1 = 0 keta = 0.102921143491894
+ lketa = -2.27421572219952E-7 wketa = -4.148835871890074E-7 pketa = 7.652982937119822E-13
+ a1 = 0 a2 = 0.8 rdsw = 547.88
+ rdswmin = 0 rdw = 0 rdwmin = 0
+ rsw = 0 rswmin = 0 prwb = -0.32348
+ prwg = 0.1376 wr = 1 voff = -0.306431699428405
+ lvoff = 1.083682108835517E-7 wvoff = 2.119386897952568E-7 pvoff = -3.727949086955869E-13
+ voffl = 0 minv = 0 nfactor = -0.352535582831901
+ lnfactor = 2.814484419326155E-6 wnfactor = 6.47398133412741E-6 pnfactor = -9.834927092594922E-12
+ eta0 = -0.743360113731169 leta0 = 1.267879396594277E-6 weta0 = 1.19978444499777E-6
+ peta0 = -1.233364012044367E-12 etab = -34.73287845433074 letab = 7.064723501432017E-5
+ wetab = 1.731583726622347E-4 petab = -3.522119700400089E-10 dsub = -0.648150933534041
+ ldsub = 9.335682618617912E-7 wdsub = 4.527488580463324E-6 pdsub = -4.65420393085333E-12
+ cit = 1E-5 cdsc = 1.3E-4 cdscb = 7.8E-4
+ cdscd = 0 pclm = 1.856015056145942 lpclm = -1.791981062492511E-6
+ wpclm = -4.947898535538428E-6 ppclm = 6.664380516990764E-12 pdiblc1 = 0.391067255322459
+ lpdiblc1 = -2.16438098688308E-9 wpdiblc1 = 3.946863256680938E-8 ppdiblc1 = -8.004191322189863E-14
+ pdiblc2 = 1.080841502366062E-3 lpdiblc2 = -6.690572543342833E-10 wpdiblc2 = -3.244700149332047E-9
+ ppdiblc2 = 3.335512817111553E-15 pdiblcb = -0.121567847713041 lpdiblcb = 1.242085294348064E-7
+ wpdiblcb = 3.572138976709622E-7 ppdiblcb = -3.673223186987996E-13 drout = 0.220528215552784
+ ldrout = 6.884447051975413E-7 wdrout = 4.014750470548685E-7 pdrout = -8.141865777267086E-13
+ pscbe1 = 7.41617730058829E8 lpscbe1 = 60.01627291228452 wpscbe1 = 174.29397330066644
+ ppscbe1 = -1.791721130254055E-4 pscbe2 = 1.328113393333894E-8 lpscbe2 = -6.482982835595877E-15
+ wpscbe2 = -7.569241086328748E-15 ppscbe2 = 8.98654949167111E-21 pvag = 0
+ delta = 0.01 fprout = 0 pdits = 0
+ pditsl = 0 pditsd = 0 lambda = 0
+ vtl = 0 lc = 5E-9 xn = 3
+ alpha0 = 2.500480180437411E-10 lalpha0 = -1.542475619727493E-16 walpha0 = -7.48048218780726E-16
+ palpha0 = 7.68984592327961E-22 alpha1 = 1E-10 beta0 = 12.627459192695833
+ lbeta0 = -3.718261244461256E-6 wbeta0 = -2.548647990510634E-5 pbeta0 = 2.579055743822103E-11
+ aigbacc = 0.43 bigbacc = 0.054 cigbacc = 0.075
+ nigbacc = 1 aigbinv = 0.35 bigbinv = 0.03
+ cigbinv = 6E-3 eigbinv = 1.1 nigbinv = 3
+ aigc = 0.43 bigc = 0.054 cigc = 0.075
+ aigsd = 0.43 bigsd = 0.054 cigsd = 0.075
+ dlcig = 0 nigc = 1 poxedge = 1
+ pigcd = 1 ntox = 1 toxref = 4.23E-9
+ agidl = -7.833916881047184E-11 lagidl = 1.833305254671393E-16 wagidl = 8.890907011422095E-16
+ pagidl = -9.139745716857775E-22 bgidl = 2.579670906362648E9 lbgidl = -1.458385786956723E3
+ wbgidl = -5.324886023134673E3 pbgidl = 5.588794453990953E-3 cgidl = 300
+ egidl = 0.1 noia = 1.5E42 noib = 0
+ noic = 0 em = 4.1E7 af = 1
+ ef = 1 kf = 0 lintnoi = -2E-7
+ tnoia = 2.5E7 tnoib = 0 ntnoi = 1
+ rnoia = 0.69 rnoib = 0.34 xpart = 0
+ cgso = {5.248925E-11/sw_func_tox_lv_ratio} cgdo = {5.248925E-11/sw_func_tox_lv_ratio} cgbo = {0/sw_func_tox_lv_ratio}
+ ckappas = 0.6 cf = 1.2E-11 clc = 1E-7
+ cle = 0.6 dlc = -3E-9 dwc = 0
+ vfbcv = -0.14469 noff = 3.9 voffcv = -0.10701
+ acde = 0.8 moin = 18.13 cgsl = {9.548271750000001E-12/sw_func_tox_lv_ratio}
+ cgdl = {9.548271750000001E-12/sw_func_tox_lv_ratio} ijthsrev = 0.1 ijthsfwd = 0.1
+ xjbvs = 1 bvs = 12.69 jss = 2.1483E-5
+ jsws = 8.040000000000001E-10 cjs = {sw_psd_nw_cj} mjs = 0.34629
+ mjsws = 0.29781 cjsws = {9.888891999999999E-11*sw_func_psd_nw_cj} cjswgs = {2.39155046E-10*sw_func_psd_nw_cj}
+ mjswgs = 0.9274 pbs = 0.6587 pbsws = 0.7418
+ pbswgs = 1.4338 xrcrg1 = 12 xrcrg2 = 1
+ rbpb = 50 rbpd = 50 rbps = 50
+ rbdb = 50 rbsb = 50 gbmin = 1E-12
+ tnom = 30 ute = 1.670237768303806 lute = -1.707494838652118E-6
+ wute = -1.007721252351072E-5 pute = 9.082322303899036E-12 kt1 = -0.390580576897025
+ lkt1 = -1.232424173078632E-7 wkt1 = -3.277669339627362E-7 pkt1 = 5.237706131868346E-13
+ kt1l = 0 kt2 = -0.011103859332743 lkt2 = -3.382303090869067E-8
+ wkt2 = -1.530647498158349E-7 pkt2 = 1.383550858601101E-13 ua1 = 3.618523894906307E-9
+ lua1 = 7.741202188209199E-16 wua1 = -1.264138616422565E-14 pua1 = 3.529779289185387E-22
+ ub1 = -6.778809423915077E-19 lub1 = -3.260151616121557E-24 wub1 = 4.172385560816075E-24
+ pub1 = 9.096946743490563E-30 uc1 = 7.196925332990231E-10 luc1 = -9.134512205846606E-16
+ wuc1 = -2.377290250098017E-15 puc1 = 3.252030268119758E-21 at = 3.539837924110048E5
+ lat = -0.398186471824882 wat = -1.090791310109455 pat = 1.422551846420603E-6
+ prt = 0 njs = 1.3632 xtis = 5.2
+ tpb = 2.0386E-3 tpbsw = 1.246E-3 tpbswg = 0
+ tcj = 1.2407E-3 tcjsw = 3.7357E-4 tcjswg = 2E-12
+ tvoff = 0 tvfbsdoff = 0 saref = 3E-6
+ sbref = 3E-6 wlod = 0 ku0 = 4.5E-8
+ kvsat = 0.5 kvth0 = 3.29E-8 tku0 = 0
+ llodku0 = 0 wlodku0 = 1 llodvth = 0
+ wlodvth = 1 lku0 = 0 wku0 = 2.5E-7
+ pku0 = 0 lkvth0 = 0 wkvth0 = 2E-7
+ pkvth0 = 0 stk2 = 0 lodk2 = 1
+ steta0 = 0 lodeta0 = 1

.model pshort_model.21 pmos
+ level = 54 lmin = 5E-7 lmax = 1E-6 wmin = 3E-6
+ wmax = 5E-6 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 4.23E-9
+ toxm = 4.23E-9 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 9.999999999999999E22 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {7.3039E-9+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {-1.3994E-8-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = -5.722E-9 dwb = -1.7864E-8 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = -1.093165510714208 lvth0 = 4.442651674247551E-8
+ wvth0 = 1.602593179624926E-7 pvth0 = -5.482247955003356E-14 k1 = 0.607856353255918
+ lk1 = -4.246813621917696E-8 wk1 = -2.84503246138047E-7 pk1 = 2.925895888611626E-14
+ k2 = -0.050323199602866 lk2 = 2.13660121821936E-8 wk2 = 1.072155717306086E-7
+ pk2 = -1.464552429812082E-14 k3 = -15.845 k3b = 2
+ w0 = 0 lpe0 = 0 lpeb = 0
+ vbm = -3 dvtp0 = 0 dvtp1 = 0
+ dvt0 = 4.4955 dvt1 = 0.294 dvt2 = 0.015
+ dvt0w = -4.9772 dvt1w = 1.1472E6 dvt2w = -8.96E-3
+ vfbsdoff = 0 u0 = 0.013462610976617 lu0 = -3.723808244630017E-9
+ wu0 = -2.168249342012874E-8 pu0 = 1.248286815729529E-14 ua = 3.946086109004071E-11
+ lua = -8.590723847503741E-16 wua = -4.630517495500919E-15 pua = 3.038622991504178E-21
+ ub = 6.115802936477759E-19 lub = 4.859652236346731E-25 wub = 2.547810935883782E-24
+ pub = -1.741254283956528E-30 uc = -4.250316955442275E-11 luc = 1.242180552153126E-17
+ wuc = -3.528268147830322E-17 puc = 3.72598476010526E-23 ud = 0
+ up = 0 lp = 1 eu = 1.67
+ vsat = -1.710667501657778E5 lvsat = 0.126608240241404 wvsat = 0.710907771934883
+ pvsat = -3.419800101070378E-7 a0 = -0.457754550615158 la0 = 6.370994897384339E-7
+ wa0 = 4.652882874594223E-6 pa0 = -2.052831846420689E-12 ags = 3.241219642825108
+ lags = -1.334857542523166E-6 wags = -8.90585793571434E-6 pags = 5.158593613831072E-12
+ b0 = 0 b1 = 0 keta = -0.226023486691235
+ lketa = 1.107295602727426E-7 wketa = 6.652891028508006E-7 pketa = -3.451062695766599E-13
+ a1 = 0 a2 = 0.858265210704412 la2 = -5.989593742160744E-8
+ wa2 = -3.03802735891508E-7 pa2 = 3.123055668636395E-13 rdsw = 547.88
+ rdswmin = 0 rdw = 0 rdwmin = 0
+ rsw = 0 rswmin = 0 prwb = -0.32348
+ prwg = 0.1376 wr = 1 voff = -0.187819540799715
+ lvoff = -1.356366484083803E-8 wvoff = -1.762617072360474E-7 pvoff = 2.627044104782963E-14
+ voffl = 0 minv = 0 nfactor = 2.937207499694352
+ lnfactor = -5.673319925938434E-7 wnfactor = -5.277388633760581E-6 pnfactor = 2.245340217954319E-12
+ eta0 = 0.49 etab = 69.88385339188537 letab = -3.689750992280787E-5
+ wetab = -3.484110660806274E-4 petab = 1.839551541543885E-10 dsub = 0.222046819523637
+ ldsub = 3.901541409153499E-8 wdsub = 2.085228671296553E-8 pdsub = -2.143590051348801E-14
+ cit = 1E-5 cdsc = 1.3E-4 cdscb = 7.8E-4
+ cdscd = 0 pclm = -0.428421300191785 lpclm = 5.563920985863959E-7
+ wpclm = 3.163984906968423E-6 ppclm = -1.674538319304969E-12 pdiblc1 = 1.046479857946062
+ lpdiblc1 = -6.759206715327156E-7 wpdiblc1 = -1.41190780375686E-6 ppdiblc1 = 1.411955646801597E-12
+ pdiblc2 = 6.781238892525484E-4 lpdiblc2 = -2.550683806649488E-10 wpdiblc2 = -1.236994902113319E-9
+ ppdiblc2 = 1.271615915433667E-15 pdiblcb = 0.236071081599945 lpdiblcb = -2.434399982317916E-7
+ wpdiblcb = -2.214369196451319E-10 ppdiblcb = 1.169160363295939E-16 drout = 0.774314128894433
+ ldrout = 1.191594317132862E-7 wdrout = -8.029500941097368E-7 pdrout = 4.239480142888117E-13
+ pscbe1 = 8E8 pscbe2 = 2.64032820157266E-8 lpscbe2 = -1.99723935985134E-14
+ wpscbe2 = -6.299508687837984E-14 ppscbe2 = 6.596365385575012E-20 pvag = 0
+ delta = 0.01 fprout = 0 pdits = 0
+ pditsl = 0 pditsd = 0 lambda = 0
+ vtl = 0 lc = 5E-9 xn = 3
+ alpha0 = 1E-10 alpha1 = 1E-10 beta0 = 8.540898913636909
+ lbeta0 = 4.826736836879706E-7 wbeta0 = -6.013005679619147E-7 pbeta0 = 2.088917017886097E-13
+ aigbacc = 0.43 bigbacc = 0.054 cigbacc = 0.075
+ nigbacc = 1 aigbinv = 0.35 bigbinv = 0.03
+ cigbinv = 6E-3 eigbinv = 1.1 nigbinv = 3
+ aigc = 0.43 bigc = 0.054 cigc = 0.075
+ aigsd = 0.43 bigsd = 0.054 cigsd = 0.075
+ dlcig = 0 nigc = 1 poxedge = 1
+ pigcd = 1 ntox = 1 toxref = 4.23E-9
+ agidl = 2.695399931777061E-10 lagidl = -1.742850785067638E-16 wagidl = -8.452233595761894E-16
+ pagidl = 8.688794709640077E-22 bgidl = 7.535211413764509E8 lbgidl = 418.87425765190875
+ wbgidl = 1.95373370342503E3 pbgidl = -1.893539281475704E-3 cgidl = 300
+ egidl = 0.1 noia = 1.5E42 noib = 0
+ noic = 0 em = 4.1E7 af = 1
+ ef = 1 kf = 0 lintnoi = -2E-7
+ tnoia = 2.5E7 tnoib = 0 ntnoi = 1
+ rnoia = 0.69 rnoib = 0.34 xpart = 0
+ cgso = {5.248925E-11/sw_func_tox_lv_ratio} cgdo = {5.248925E-11/sw_func_tox_lv_ratio} cgbo = {0/sw_func_tox_lv_ratio}
+ ckappas = 0.6 cf = 1.2E-11 clc = 1E-7
+ cle = 0.6 dlc = -3E-9 dwc = 0
+ vfbcv = -0.14469 noff = 3.9 voffcv = -0.10701
+ acde = 0.8 moin = 18.13 cgsl = {9.548271750000001E-12/sw_func_tox_lv_ratio}
+ cgdl = {9.548271750000001E-12/sw_func_tox_lv_ratio} ijthsrev = 0.1 ijthsfwd = 0.1
+ xjbvs = 1 bvs = 12.69 jss = 2.1483E-5
+ jsws = 8.040000000000001E-10 cjs = {sw_psd_nw_cj} mjs = 0.34629
+ mjsws = 0.29781 cjsws = {9.888891999999999E-11*sw_func_psd_nw_cj} cjswgs = {2.39155046E-10*sw_func_psd_nw_cj}
+ mjswgs = 0.9274 pbs = 0.6587 pbsws = 0.7418
+ pbswgs = 1.4338 xrcrg1 = 12 xrcrg2 = 1
+ rbpb = 50 rbpd = 50 rbps = 50
+ rbdb = 50 rbsb = 50 gbmin = 1E-12
+ tnom = 30 ute = 0.35438874550195 lute = -3.548178334000834E-7
+ wute = -2.5538624874394E-6 pute = 1.348408747018154E-12 kt1 = -0.512587569822165
+ lkt1 = 2.1793073352651E-9 wkt1 = 3.736602765526986E-7 pkt1 = -1.972881420965062E-13
+ kt1l = 0 kt2 = -0.032198126624877 lkt2 = -1.213837726358451E-8
+ wkt2 = -3.798728034714076E-8 pkt2 = 2.005682817592615E-14 ua1 = 8.693303270092573E-9
+ lua1 = -4.44269208151806E-15 wua1 = -2.615858028798673E-14 pua1 = 1.424849128181544E-20
+ ub1 = -8.433199018545431E-18 lub1 = 4.712222302347765E-24 wub1 = 2.700647192056918E-23
+ pub1 = -1.437622002529932E-29 uc1 = -3.729132016473284E-10 luc1 = 2.097343636713696E-16
+ wuc1 = 1.616408837003996E-15 puc1 = -8.534444690320656E-22 at = -1.387095871730762E5
+ lat = 0.108296410066998 wat = 0.578888246083538 pat = -2.938587011911184E-7
+ prt = 0 njs = 1.3632 xtis = 5.2
+ tpb = 2.0386E-3 tpbsw = 1.246E-3 tpbswg = 0
+ tcj = 1.2407E-3 tcjsw = 3.7357E-4 tcjswg = 2E-12
+ tvoff = 0 tvfbsdoff = 0 saref = 2.75E-6
+ sbref = 2.74E-6 wlod = 0 ku0 = 4.5E-8
+ kvsat = 0.5 kvth0 = 3.29E-8 tku0 = 0
+ llodku0 = 0 wlodku0 = 1 llodvth = 0
+ wlodvth = 1 lku0 = 0 wku0 = 2.5E-7
+ pku0 = 0 lkvth0 = 0 wkvth0 = 2E-7
+ pkvth0 = 0 stk2 = 0 lodk2 = 1
+ steta0 = 0 lodeta0 = 1

.model pshort_model.22 pmos
+ level = 54 lmin = 2.5E-7 lmax = 5E-7 wmin = 3E-6
+ wmax = 5E-6 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 4.23E-9
+ toxm = 4.23E-9 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 9.999999999999999E22 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {7.3039E-9+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {-1.3994E-8-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = -5.722E-9 dwb = -1.7864E-8 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = -1.003336200261516 lvth0 = -3.002281224820515E-9
+ wvth0 = 1.181299598959398E-8 pvth0 = 2.355539709579281E-14 k1 = 0.111235728789203
+ lk1 = 2.19741594051755E-7 wk1 = -4.913825247517912E-8 pk1 = -9.501093338795401E-14
+ k2 = 0.127938719360873 lk2 = -7.275414188763273E-8 wk2 = 2.343740963099267E-8
+ pk2 = 2.958833995253117E-14 k3 = -15.845 k3b = 2
+ w0 = 0 lpe0 = 0 lpeb = 0
+ vbm = -3 dvtp0 = 0 dvtp1 = 0
+ dvt0 = 4.4955 dvt1 = 0.294 dvt2 = 0.015
+ dvt0w = -4.9772 dvt1w = 1.1472E6 dvt2w = -8.96E-3
+ vfbsdoff = 0 u0 = 8.735545691710372E-3 lu0 = -1.227974498982525E-9
+ wu0 = 4.12146199148249E-9 pu0 = -1.141310652570495E-15 ua = -9.35894198245188E-10
+ lua = -3.440966176820854E-16 wua = 1.669498665019787E-15 pua = -2.877099410568281E-22
+ ub = 1.02366082295916E-18 lub = 2.683916491246139E-25 wub = -9.77010244914082E-25
+ pub = 1.198090016505741E-31 uc = -5.108559730520197E-11 luc = 1.695322438480968E-17
+ wuc = 1.287446032330907E-16 puc = -4.934459039914687E-23 ud = 0
+ up = 0 lp = 1 eu = 1.67
+ vsat = 1.350821712071161E5 lvsat = -0.035034716456427 wvsat = -0.282665037304663
+ pvsat = 1.826145102977316E-7 a0 = 0.559400242467097 la0 = 1.000539648485201E-7
+ wa0 = 3.004304171215358E-6 pa0 = -1.182402073981089E-12 ags = -3.265263624877713
+ lags = 2.100487545024711E-6 wags = 1.306641489221675E-5 pags = -6.442502772042607E-12
+ b0 = 0 b1 = 0 keta = 0.117680960981484
+ lketa = -7.074226364508113E-8 wketa = -1.735940961075201E-7 pketa = 9.781399287494585E-14
+ a1 = 0 a2 = 0.683469578591175 la2 = 3.239405878659638E-8
+ wa2 = 6.076054717830163E-7 pa2 = -1.689070298900171E-13 rdsw = 547.88
+ rdswmin = 0 rdw = 0 rdwmin = 0
+ rsw = 0 rswmin = 0 prwb = -0.32348
+ prwg = 0.1376 wr = 1 voff = -0.205339729331252
+ lvoff = -4.313215538448761E-9 wvoff = -2.008550334856293E-8 pvoff = -5.61887204903155E-14
+ voffl = 0 minv = 0 nfactor = 1.385008848530791
+ lnfactor = 2.522102688367026E-7 wnfactor = -6.039568290103188E-7 pnfactor = -2.221756937721624E-13
+ eta0 = 0.353485933730394 leta0 = 7.207778882155675E-8 weta0 = 1.061878373704399E-6
+ peta0 = -5.606590387754383E-13 etab = 5.142315273416213E-3 letab = -2.389018889667685E-9
+ wetab = -1.812337018332253E-8 petab = 7.861118586549685E-15 dsub = 0.290725058975033
+ ldsub = 2.754127800071418E-9 wdsub = -7.097589907723811E-7 pdsub = 3.643180866634452E-13
+ cit = 1E-5 cdsc = 1.3E-4 cdscb = 7.8E-4
+ cdscd = 0 pclm = 0.812502089886036 lpclm = -9.880056029401221E-8
+ wpclm = -1.317197402704583E-6 ppclm = 6.914721660146625E-13 pdiblc1 = -0.87109547305574
+ lpdiblc1 = 3.365360923322638E-7 wpdiblc1 = 2.507697380675921E-6 ppdiblc1 = -6.575488553166974E-13
+ pdiblc2 = -5.00165762792038E-3 lpdiblc2 = 2.743788103024151E-9 wpdiblc2 = -7.154077808046222E-9
+ ppdiblc2 = 4.395764684771368E-15 pdiblcb = -0.612965135720229 lpdiblcb = 2.04840936078652E-7
+ wpdiblcb = 8.25454995976688E-7 ppdiblcb = -4.358303324157395E-13 drout = 1.010833016324188
+ ldrout = -5.719702622975275E-9 wdrout = 1.342271233284695E-6 pdrout = -7.087031039195196E-13
+ pscbe1 = 8E8 pscbe2 = -4.685776953334532E-8 lpscbe2 = 1.870856248677798E-14
+ wpscbe2 = 1.680434990578746E-13 ppscbe2 = -5.602194705556099E-20 pvag = 0
+ delta = 0.01 fprout = 0 pdits = 0
+ pditsl = 0 pditsd = 0 lambda = 0
+ vtl = 0 lc = 5E-9 xn = 3
+ alpha0 = -2.32128195859522E-8 lalpha0 = 1.230888898754773E-14 walpha0 = 6.959790975190892E-14
+ palpha0 = -3.674686117409088E-20 alpha1 = 3.771758413787202E-10 lalpha1 = -1.463455181378677E-16
+ walpha1 = -8.274785948804684E-16 palpha1 = 4.368987683537487E-22 beta0 = -8.501510078309245
+ lbeta0 = 9.480861122527635E-6 wbeta0 = 5.494065380089383E-5 pbeta0 = -2.911659370151479E-11
+ aigbacc = 0.43 bigbacc = 0.054 cigbacc = 0.075
+ nigbacc = 1 aigbinv = 0.35 bigbinv = 0.03
+ cigbinv = 6E-3 eigbinv = 1.1 nigbinv = 3
+ aigc = 0.43 bigc = 0.054 cigc = 0.075
+ aigsd = 0.43 bigsd = 0.054 cigsd = 0.075
+ dlcig = 0 nigc = 1 poxedge = 1
+ pigcd = 1 ntox = 1 toxref = 4.23E-9
+ agidl = 3.848841627980795E-9 lagidl = -2.064113390063176E-15 wagidl = -1.868944581117075E-14
+ pagidl = 1.029041479473652E-20 bgidl = 3.475238682106924E7 lbgidl = 798.3755348320954
+ wbgidl = 2.881642695452997E3 pbgidl = -2.383464094358566E-3 cgidl = 626.2555741959075
+ lcgidl = -1.722590281085488E-4 wcgidl = -1.798780830597812E-4 pcgidl = 9.497346931856777E-11
+ egidl = 2.201119726620335 legidl = -1.109366002218817E-6 wegidl = -1.047490589635915E-5
+ pegidl = 5.530624614406873E-12 noia = 1.5E42 noib = 0
+ noic = 0 em = 4.1E7 af = 1
+ ef = 1 kf = 0 lintnoi = -2E-7
+ tnoia = 2.5E7 tnoib = 0 ntnoi = 1
+ rnoia = 0.69 rnoib = 0.34 xpart = 0
+ cgso = {5.248925E-11/sw_func_tox_lv_ratio} cgdo = {5.248925E-11/sw_func_tox_lv_ratio} cgbo = {0/sw_func_tox_lv_ratio}
+ ckappas = 0.6 cf = 1.2E-11 clc = 1E-7
+ cle = 0.6 dlc = -3E-9 dwc = 0
+ vfbcv = -0.14469 noff = 3.9 voffcv = -0.10701
+ acde = 0.8 moin = 18.13 cgsl = {9.548271750000001E-12/sw_func_tox_lv_ratio}
+ cgdl = {9.548271750000001E-12/sw_func_tox_lv_ratio} ijthsrev = 0.1 ijthsfwd = 0.1
+ xjbvs = 1 bvs = 12.69 jss = 2.1483E-5
+ jsws = 8.040000000000001E-10 cjs = {sw_psd_nw_cj} mjs = 0.34629
+ mjsws = 0.29781 cjsws = {9.888891999999999E-11*sw_func_psd_nw_cj} cjswgs = {2.39155046E-10*sw_func_psd_nw_cj}
+ mjswgs = 0.9274 pbs = 0.6587 pbsws = 0.7418
+ pbswgs = 1.4338 xrcrg1 = 12 xrcrg2 = 1
+ rbpb = 50 rbpd = 50 rbps = 50
+ rbdb = 50 rbsb = 50 gbmin = 1E-12
+ tnom = 30 ute = -0.33723371376 lute = 1.03505256207149E-8
+ kt1 = -0.386136323069855 lkt1 = -6.458543353499341E-8 wkt1 = -2.797705129290854E-7
+ pkt1 = 1.47715473580402E-13 kt1l = 0 kt2 = 0.11033875387042
+ lkt2 = -8.739613972253508E-8 wkt2 = -4.753533536150338E-7 pkt2 = 2.509808664684945E-13
+ ua1 = 4.578041050702511E-10 lua1 = -9.444734837625375E-17 wua1 = 1.469852623710351E-15
+ pua1 = -3.389897543656737E-22 ub1 = 5.581698006953996E-19 lub1 = -3.51125377855635E-26
+ wub1 = -3.385108283516156E-25 pub1 = 6.16027263378785E-32 uc1 = 1.052515366186829E-11
+ luc1 = 7.28351332837748E-18 wuc1 = 1.199227491023493E-16 puc1 = -6.33177724530512E-23
+ at = 6.722820410397112E4 lat = -4.362724737879052E-4 wat = 0.078519097860064
+ pat = -2.966979535890307E-8 prt = 0 njs = 1.3632
+ xtis = 5.2 tpb = 2.0386E-3 tpbsw = 1.246E-3
+ tpbswg = 0 tcj = 1.2407E-3 tcjsw = 3.7357E-4
+ tcjswg = 2E-12 tvoff = 0 tvfbsdoff = 0
+ saref = 1.75E-6 sbref = 1.74E-6 wlod = 0
+ ku0 = 4.5E-8 kvsat = 0.5 kvth0 = 3.29E-8
+ tku0 = 0 llodku0 = 0 wlodku0 = 1
+ llodvth = 0 wlodvth = 1 lku0 = 0
+ wku0 = 2.5E-7 pku0 = 0 lkvth0 = 0
+ wkvth0 = 2E-7 pkvth0 = 0 stk2 = 0
+ lodk2 = 1 steta0 = 0 lodeta0 = 1

.model pshort_model.23 pmos
+ level = 54 lmin = 1.8E-7 lmax = 2.5E-7 wmin = 3E-6
+ wmax = 5E-6 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 4.23E-9
+ toxm = 4.23E-9 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 9.999999999999999E22 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {7.3039E-9+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {-1.3994E-8-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = -5.722E-9 dwb = -1.7864E-8 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = -0.948983603979548 lvth0 = -1.811165076005212E-8
+ wvth0 = 1.497764246363518E-7 pvth0 = -1.47967805068621E-14 k1 = 0.517108815050108
+ lk1 = 1.069137465482586E-7 wk1 = -1.610315571141452E-6 pk1 = 3.38977627073446E-13
+ k2 = 9.897414527498621E-3 lk2 = -3.994007563961272E-8 wk2 = 5.759450910010071E-7
+ pk2 = -1.240021653761564E-13 k3 = -15.845 k3b = 2
+ w0 = 0 lpe0 = 0 lpeb = 0
+ vbm = -3 dvtp0 = 0 dvtp1 = 0
+ dvt0 = 4.4955 dvt1 = 0.294 dvt2 = 0.015
+ dvt0w = -4.9772 dvt1w = 1.1472E6 dvt2w = -8.96E-3
+ vfbsdoff = 0 u0 = 6.425365683448595E-3 lu0 = -5.857721788458498E-10
+ wu0 = 5.902979642914947E-10 pu0 = -1.596894269797248E-16 ua = -1.768314166309505E-9
+ lua = -1.12693855599822E-16 wua = 1.899142900817894E-15 pua = -3.515482828778722E-22
+ ub = 1.86129873909603E-18 lub = 3.553836009355797E-26 wub = -2.310525467047572E-24
+ pub = 4.905102312210186E-31 uc = 3.880909642344183E-11 luc = -8.036421735428552E-18
+ wuc = -1.943732216979982E-16 puc = 4.047828751779668E-23 ud = 0
+ up = 0 lp = 1 eu = 1.67
+ vsat = -2.197988870015829E5 lvsat = 0.063617959152893 wvsat = 1.389120025142025
+ pvsat = -2.821216756416984E-7 a0 = 3.755546059110616 la0 = -7.884362184285784E-7
+ wa0 = -1.317554247407782E-5 pa0 = 3.31540113525067E-12 ags = 13.325692006745781
+ lags = -2.511599029099041E-6 wags = -4.014566041407223E-5 pags = 8.349815618202055E-12
+ b0 = 0 b1 = -1.560790734647861E-23 lb1 = 4.338810947432896E-30
+ wb1 = 4.659572485049995E-29 pb1 = -1.295305235974078E-35 keta = -0.073204668515808
+ lketa = -1.767834927238786E-8 wketa = -9.073094438554571E-7 pketa = 3.017780549646994E-13
+ a1 = 0 a2 = 0.518565270761412 la2 = 7.823547751157656E-8
+ wa2 = 1.976692699697488E-6 pa2 = -5.494968502035054E-13 rdsw = 547.88
+ rdswmin = 0 rdw = 0 rdwmin = 0
+ rsw = 0 rswmin = 0 prwb = -0.32348
+ prwg = 0.1376 wr = 1 voff = 0.095759986126976
+ lvoff = -8.80153232392507E-8 wvoff = -7.04408829512716E-7 pvoff = 1.34044952303405E-13
+ voffl = 0 minv = 0 nfactor = 2.171126613065283
+ lnfactor = 3.367896370928842E-8 wnfactor = -3.366560078548638E-6 pnfactor = 5.457948583604958E-13
+ eta0 = 1.776509391992726 leta0 = -3.235056562938724E-7 weta0 = -3.445665607346728E-6
+ peta0 = 6.923840974290025E-13 etab = 0.051845539421046 letab = -1.537195476401896E-8
+ wetab = 5.396563220249986E-7 petab = -1.471949424910571E-13 dsub = 0.153984768260276
+ ldsub = 4.076628773528526E-8 wdsub = 3.08029943039803E-6 pdsub = -6.892726737208749E-13
+ cit = 1E-5 cdsc = 1.3E-4 cdscb = 7.8E-4
+ cdscd = 0 pclm = -0.109830324704987 lpclm = 1.575967829733171E-7
+ wpclm = 4.798045881657205E-6 ppclm = -1.008492084118502E-12 pdiblc1 = 0.737367328973287
+ lpdiblc1 = -1.105972650781813E-7 wpdiblc1 = 7.852997907286824E-7 ppdiblc1 = -1.787429940824446E-13
+ pdiblc2 = 5.948617714430884E-3 lpdiblc2 = -3.002570388453927E-10 wpdiblc2 = 3.86282018634308E-8
+ ppdiblc2 = -8.331159676543187E-15 pdiblcb = 1.046682042566234 lpdiblcb = -2.565210637188449E-7
+ wpdiblcb = -4.602111186680052E-6 ppdiblcb = 1.072967935568642E-12 drout = 1.617856330075446
+ ldrout = -1.7446489956606E-7 wdrout = -6.753872167532854E-6 pdrout = 1.541927607786949E-12
+ pscbe1 = 8E8 pscbe2 = 5.385798880490326E-8 lpscbe2 = -9.289209742155073E-15
+ wpscbe2 = -1.354639777504796E-13 ppscbe2 = 2.834948940743981E-20 pvag = 0
+ delta = 0.01 fprout = 0 pdits = 0
+ pditsl = 0 pditsd = 0 lambda = 0
+ vtl = 0 lc = 5E-9 xn = 3
+ alpha0 = 8.336006994982924E-8 lalpha0 = -1.731709542872508E-14 walpha0 = -2.485639633996746E-13
+ palpha0 = 5.169832161957153E-20 alpha1 = -8.899137192097142E-10 lalpha1 = 2.058901746309901E-16
+ walpha1 = 2.955280696001672E-15 palpha1 = -6.146629213999957E-22 beta0 = 76.16501835810192
+ lbeta0 = -1.405541778445343E-5 wbeta0 = -1.977116041345593E-4 pbeta0 = 4.111770217744595E-11
+ aigbacc = 0.43 bigbacc = 0.054 cigbacc = 0.075
+ nigbacc = 1 aigbinv = 0.35 bigbinv = 0.03
+ cigbinv = 6E-3 eigbinv = 1.1 nigbinv = 3
+ aigc = 0.43 bigc = 0.054 cigc = 0.075
+ aigsd = 0.43 bigsd = 0.054 cigsd = 0.075
+ dlcig = 0 nigc = 1 poxedge = 1
+ pigcd = 1 ntox = 1 toxref = 4.23E-9
+ agidl = -1.360571860329356E-8 lagidl = 2.788044899508319E-15 wagidl = 6.832838262025462E-14
+ pagidl = -1.389949729525856E-20 bgidl = 7.882249052550169E9 lbgidl = -1.383134368280606E3
+ wbgidl = -2.054621263994066E4 pbgidl = 4.129198554616847E-3 cgidl = -865.1984792710978
+ lcgidl = 2.423473013066371E-4 wcgidl = 6.424217252135043E-4 pcgidl = -1.336160097837063E-10
+ egidl = -7.403999023644049 legidl = 1.560741748929678E-6 wegidl = 3.741037820128266E-5
+ pegidl = -7.780909741328378E-12 noia = 1.5E42 noib = 0
+ noic = 0 em = 4.1E7 af = 1
+ ef = 1 kf = 0 lintnoi = -2E-7
+ tnoia = 2.5E7 tnoib = 0 ntnoi = 1
+ rnoia = 0.69 rnoib = 0.34 xpart = 0
+ cgso = {5.248925E-11/sw_func_tox_lv_ratio} cgdo = {5.248925E-11/sw_func_tox_lv_ratio} cgbo = {0/sw_func_tox_lv_ratio}
+ ckappas = 0.6 cf = 1.2E-11 clc = 1E-7
+ cle = 0.6 dlc = -3E-9 dwc = 0
+ vfbcv = -0.14469 noff = 3.9 voffcv = -0.10701
+ acde = 0.8 moin = 18.13 cgsl = {9.548271750000001E-12/sw_func_tox_lv_ratio}
+ cgdl = {9.548271750000001E-12/sw_func_tox_lv_ratio} ijthsrev = 0.1 ijthsfwd = 0.1
+ xjbvs = 1 bvs = 12.69 jss = 2.1483E-5
+ jsws = 8.040000000000001E-10 cjs = {sw_psd_nw_cj} mjs = 0.34629
+ mjsws = 0.29781 cjsws = {9.888891999999999E-11*sw_func_psd_nw_cj} cjswgs = {2.39155046E-10*sw_func_psd_nw_cj}
+ mjswgs = 0.9274 pbs = 0.6587 pbsws = 0.7418
+ pbswgs = 1.4338 xrcrg1 = 12 xrcrg2 = 1
+ rbpb = 50 rbpd = 50 rbps = 50
+ rbdb = 50 rbsb = 50 gbmin = 1E-12
+ tnom = 30 ute = -0.3 kt1 = -0.901477142942004
+ lkt1 = 7.86731302996255E-8 wkt1 = 1.662514347301351E-6 pkt1 = -3.922164101453367E-13
+ kt1l = 0 kt2 = -0.47506577056286 lkt2 = 7.533929321562332E-8
+ wkt2 = 1.778617289791069E-6 pkt2 = -3.755959247506813E-13 ua1 = 6.881935177164556E-11
+ lua1 = 1.368574522371898E-17 wua1 = 9.944519542045618E-16 pua1 = -2.068340730510984E-22
+ ub1 = 5.482154452878463E-19 lub1 = -3.234534643452858E-26 wub1 = -4.642745973418632E-25
+ pub1 = 9.656354495193943E-32 uc1 = 3.672597286405501E-11 wuc1 = -1.078488541792715E-16
+ at = 1.694275599550746E5 lat = -0.028846467008124 wat = -0.445404220299908
+ pat = 1.159746000097512E-7 prt = 0 njs = 1.3632
+ xtis = 5.2 tpb = 2.0386E-3 tpbsw = 1.246E-3
+ tpbswg = 0 tcj = 1.2407E-3 tcjsw = 3.7357E-4
+ tcjswg = 2E-12 tvoff = 0 tvfbsdoff = 0
+ saref = 1.25E-6 sbref = 1.24E-6 wlod = 0
+ ku0 = 4.5E-8 kvsat = 0.5 kvth0 = 3.29E-8
+ tku0 = 0 llodku0 = 0 wlodku0 = 1
+ llodvth = 0 wlodvth = 1 lku0 = 0
+ wku0 = 2.5E-7 pku0 = 0 lkvth0 = 0
+ wkvth0 = 2E-7 pkvth0 = 0 stk2 = 0
+ lodk2 = 1 steta0 = 0 lodeta0 = 1

.model pshort_model.24 pmos
+ level = 54 lmin = 1.5E-7 lmax = 1.8E-7 wmin = 3E-6
+ wmax = 5E-6 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 4.23E-9
+ toxm = 4.23E-9 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 9.999999999999999E22 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {7.3039E-9+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {-1.3994E-8-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = -5.722E-9 dwb = -1.7864E-8 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = -0.956083599107521 lvth0 = -1.663493697337535E-8
+ wvth0 = 4.73242028690363E-7 pvth0 = -8.207374456284779E-14 k1 = -0.296887372665633
+ lk1 = 2.7621518563888E-7 wk1 = -9.609112435829802E-7 pk1 = 2.039093197932145E-13
+ k2 = 0.396688359746296 lk2 = -1.203879507537799E-7 wk2 = 2.883206204214418E-7
+ pk2 = -6.417972698925379E-14 k3 = -15.845 k3b = 2
+ w0 = 0 lpe0 = 0 lpeb = 0
+ vbm = -3 dvtp0 = 0 dvtp1 = 0
+ dvt0 = 4.4955 dvt1 = 0.294 dvt2 = 0.015
+ dvt0w = -4.9772 dvt1w = 1.1472E6 dvt2w = -8.96E-3
+ vfbsdoff = 0 u0 = 6.724192038512655E-3 lu0 = -6.479244747829139E-10
+ wu0 = -1.148805181590539E-9 pu0 = 2.020231581259883E-16 ua = -6.946130715027984E-10
+ lua = -3.360107989064793E-16 wua = -3.328604519112609E-16 pua = 1.126816304495592E-22
+ ub = 1.256468989171684E-19 lub = 3.965331150286789E-25 wub = 1.415333929221365E-24
+ pub = -2.84423812890165E-31 uc = 8.642142495847417E-13 luc = -1.44341581852367E-19
+ wuc = -8.465162881813949E-19 puc = 2.270551130197101E-25 ud = 0
+ up = 0 lp = 1 eu = 1.67
+ vsat = 1.173347014571078E5 lvsat = -6.5017816434535E-3 wvsat = 0.67469115086003
+ pvsat = -1.335290429375348E-7 a0 = -6.860777121259114 la0 = 1.419631607210161E-6
+ wa0 = 2.386914779098207E-5 pa0 = -4.389449903598605E-12 ags = 1.25
+ b0 = 0 b1 = 3.641845047511675E-23 lb1 = -6.48204716316508E-30
+ wb1 = -1.087233579844998E-28 pb1 = 1.935145304094516E-35 keta = -0.82504886018321
+ lketa = 1.386962204641318E-7 wketa = 2.70535575118545E-6 pketa = -4.496129536214689E-13
+ a1 = 0 a2 = 2.763446467045952 la2 = -3.886728727412523E-7
+ wa2 = -1.204706080719114E-5 pa2 = 2.367275594187246E-12 rdsw = 547.88
+ rdswmin = 0 rdw = 0 rdwmin = 0
+ rsw = 0 rswmin = 0 prwb = -0.32348
+ prwg = 0.1376 wr = 1 voff = 0.079332073110952
+ lvoff = -8.459851446687401E-8 wvoff = -4.612557052930391E-7 pvoff = 8.347202030320289E-14
+ voffl = 0 minv = 0 nfactor = 3.61329944061981
+ lnfactor = -2.662756783481223E-7 wnfactor = -1.625624035294874E-5 pnfactor = 3.226693679272425E-12
+ eta0 = 0.121958650053125 leta0 = 2.062104342066128E-8 weta0 = -2.455409145336719E-6
+ peta0 = 4.864226364084649E-13 etab = -0.062358180255604 letab = 8.381048484087996E-9
+ wetab = -1.189510364452878E-6 petab = 2.124509782961036E-13 dsub = 0.883879723873454
+ ldsub = -1.110431042927883E-7 wdsub = -1.620245193041652E-6 pdsub = 2.883842014190976E-13
+ cit = 1E-5 cdsc = 1.3E-4 cdscb = 7.8E-4
+ cdscd = 0 pclm = 1.607325499451994 lpclm = -1.995510225814451E-7
+ wpclm = 4.05967044305216E-7 ppclm = -9.499239089533689E-14 pdiblc1 = 1.309850003159835
+ lpdiblc1 = -2.29666791516893E-7 wpdiblc1 = -5.136662344915637E-7 ppdiblc1 = 9.142635157106393E-14
+ pdiblc2 = 0.013260460026266 lpdiblc2 = -1.821032497599395E-9 wpdiblc2 = 3.613969838613579E-8
+ ppdiblc2 = -7.813580815307553E-15 pdiblcb = -0.185381051168264 lpdiblcb = -2.667249791943218E-10
+ wpdiblcb = 5.502928315220645E-7 ppdiblcb = 1.329728630820545E-15 drout = -0.531939906210939
+ ldrout = 2.726669200266726E-7 wdrout = 4.573441446870868E-6 pdrout = -8.14017696245652E-13
+ pscbe1 = 8E8 pscbe2 = 1.066729406212156E-8 lpscbe2 = -3.060635239933914E-16
+ wpscbe2 = -5.000543117925561E-15 ppscbe2 = 1.214660565084148E-21 pvag = 0
+ delta = 0.01 fprout = 0 pdits = 0
+ pditsl = 0 pditsd = 0 lambda = 0
+ vtl = 0 lc = 5E-9 xn = 3
+ alpha0 = 1E-10 alpha1 = 1E-10 beta0 = 11.059381197646326
+ lbeta0 = -5.142265227245942E-7 wbeta0 = 1.382518383621016E-5 pbeta0 = -2.879411279018446E-12
+ aigbacc = 0.43 bigbacc = 0.054 cigbacc = 0.075
+ nigbacc = 1 aigbinv = 0.35 bigbinv = 0.03
+ cigbinv = 6E-3 eigbinv = 1.1 nigbinv = 3
+ aigc = 0.43 bigc = 0.054 cigc = 0.075
+ aigsd = 0.43 bigsd = 0.054 cigsd = 0.075
+ dlcig = 0 nigc = 1 poxedge = 1
+ pigcd = 1 ntox = 1 toxref = 4.23E-9
+ agidl = -1.046272094996323E-9 lagidl = 1.758307391405933E-16 wagidl = 4.554872950902241E-15
+ pagidl = -6.353725661492973E-22 bgidl = 2.609694922039965E9 lbgidl = -286.5063797840492
+ wbgidl = -4.805570664637718E3 pbgidl = 8.553339114575382E-4 cgidl = 300
+ egidl = 0.1 noia = 1.5E42 noib = 0
+ noic = 0 em = 4.1E7 af = 1
+ ef = 1 kf = 0 lintnoi = -2E-7
+ tnoia = 2.5E7 tnoib = 0 ntnoi = 1
+ rnoia = 0.69 rnoib = 0.34 xpart = 0
+ cgso = {5.248925E-11/sw_func_tox_lv_ratio} cgdo = {5.248925E-11/sw_func_tox_lv_ratio} cgbo = {0/sw_func_tox_lv_ratio}
+ ckappas = 0.6 cf = 1.2E-11 clc = 1E-7
+ cle = 0.6 dlc = -3E-9 dwc = 0
+ vfbcv = -0.14469 noff = 3.9 voffcv = -0.10701
+ acde = 0.8 moin = 18.13 cgsl = {9.548271750000001E-12/sw_func_tox_lv_ratio}
+ cgdl = {9.548271750000001E-12/sw_func_tox_lv_ratio} ijthsrev = 0.1 ijthsfwd = 0.1
+ xjbvs = 1 bvs = 12.69 jss = 2.1483E-5
+ jsws = 8.040000000000001E-10 cjs = {sw_psd_nw_cj} mjs = 0.34629
+ mjsws = 0.29781 cjsws = {9.888891999999999E-11*sw_func_psd_nw_cj} cjswgs = {2.39155046E-10*sw_func_psd_nw_cj}
+ mjswgs = 0.9274 pbs = 0.6587 pbsws = 0.7418
+ pbswgs = 1.4338 xrcrg1 = 12 xrcrg2 = 1
+ rbpb = 50 rbpd = 50 rbps = 50
+ rbdb = 50 rbsb = 50 gbmin = 1E-12
+ tnom = 30 ute = -0.3 kt1 = 0.466367410217013
+ lkt1 = -2.058221226228121E-7 wkt1 = -1.459477273440099E-6 pkt1 = 2.571203830694361E-13
+ kt1l = 0 kt2 = -0.05870899307349 lkt2 = -1.125792022083558E-8
+ wkt2 = -1.888290627205475E-7 pkt2 = 3.36093072155048E-14 ua1 = 1.3462E-10
+ ub1 = 3.927E-19 uc1 = 2.925624880163569E-11 luc1 = 1.553612968294461E-18
+ wuc1 = -7.477089161012767E-16 puc1 = 1.33083214559034E-22 at = -1.237038893961348E4
+ lat = 8.965324786583927E-3 wat = 0.777862234600464 pat = -1.384501434120673E-7
+ prt = 0 njs = 1.3632 xtis = 5.2
+ tpb = 2.0386E-3 tpbsw = 1.246E-3 tpbswg = 0
+ tcj = 1.2407E-3 tcjsw = 3.7357E-4 tcjswg = 2E-12
+ tvoff = 0 tvfbsdoff = 0 saref = 1.1E-6
+ sbref = 1.1E-6 wlod = 0 ku0 = 4.5E-8
+ kvsat = 0.5 kvth0 = 3.29E-8 tku0 = 0
+ llodku0 = 0 wlodku0 = 1 llodvth = 0
+ wlodvth = 1 lku0 = 0 wku0 = 2.5E-7
+ pku0 = 0 lkvth0 = 0 wkvth0 = 2E-7
+ pkvth0 = 0 stk2 = 0 lodk2 = 1
+ steta0 = 0 lodeta0 = 1

.model pshort_model.25 pmos
+ level = 54 lmin = 8E-6 lmax = 2.02E-5 wmin = 1E-6
+ wmax = 3E-6 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 4.23E-9
+ toxm = 4.23E-9 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 9.999999999999999E22 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {7.3039E-9+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {-1.3994E-8-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = -5.722E-9 dwb = -1.7864E-8 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = -1.06157667141295 wvth0 = 4.119892409488394E-8
+ k1 = 0.389161224322262 wk1 = 1.011099069122368E-7 k2 = 0.033201497874547
+ wk2 = -3.53674454437687E-8 k3 = -15.845 k3b = 2
+ w0 = 0 lpe0 = 0 lpeb = 0
+ vbm = -3 dvtp0 = 0 dvtp1 = 0
+ dvt0 = 4.4955 dvt1 = 0.294 dvt2 = 0.015
+ dvt0w = -4.9772 dvt1w = 1.1472E6 dvt2w = -8.96E-3
+ vfbsdoff = 0 u0 = 0.014188902684328 wu0 = -7.84084208785271E-9
+ ua = 4.062596229700033E-10 wua = -1.791338295043602E-15 ub = 4.059411094322819E-19
+ wub = 9.50066767188483E-25 uc = -1.280177637498152E-10 wuc = 8.779959571155947E-17
+ ud = 0 up = 0 lp = 1
+ eu = 1.67 vsat = 5.25512371833863E4 wvsat = 2.647334795968575E-3
+ a0 = 1.058691498271 wa0 = 1.51339984652443E-7 ags = 0.129833294476556
+ wags = 1.559086312257727E-7 b0 = 0 b1 = 0
+ keta = -3.264199199107872E-3 wketa = 9.759754471616204E-9 a1 = 0
+ a2 = 0.8 rdsw = 547.88 rdswmin = 0
+ rdw = 0 rdwmin = 0 rsw = 0
+ rswmin = 0 prwb = -0.32348 prwg = 0.1376
+ wr = 1 voff = -0.25245591 voffl = 0
+ minv = 0 nfactor = 1.83670682814142 wnfactor = -2.737360685371356E-7
+ eta0 = 0.08 etab = -0.07 dsub = 0.56
+ cit = 1E-5 cdsc = 1.3E-4 cdscb = 7.8E-4
+ cdscd = 0 pclm = 0.221212410156329 wpclm = -2.162661701073159E-7
+ pdiblc1 = 0.39 pdiblc2 = 6.661719080525955E-6 wpdiblc2 = 5.529790650764066E-10
+ pdiblcb = 0.07353922 wpdiblcb = -2.94178218782084E-7 drout = 0.56
+ pscbe1 = 7.36012798315339E8 wpscbe1 = 63.037994320629814 pscbe2 = 9.430440234047E-9
+ wpscbe2 = 1.321933952830112E-15 pvag = 0 delta = 0.01
+ fprout = 0 pdits = 0 pditsl = 0
+ pditsd = 0 lambda = 0 vtl = 0
+ lc = 5E-9 xn = 3 alpha0 = 2.65936214519591E-11
+ walpha0 = -2.620514714851318E-17 alpha1 = 9.412422596166031E-17 walpha1 = -9.274927809365758E-23
+ beta0 = -0.332026142236774 wbeta0 = 2.988894197075621E-5 aigbacc = 0.43
+ bigbacc = 0.054 cigbacc = 0.075 nigbacc = 1
+ aigbinv = 0.35 bigbinv = 0.03 cigbinv = 6E-3
+ eigbinv = 1.1 nigbinv = 3 aigc = 0.43
+ bigc = 0.054 cigc = 0.075 aigsd = 0.43
+ bigsd = 0.054 cigsd = 0.075 dlcig = 0
+ nigc = 1 poxedge = 1 pigcd = 1
+ ntox = 1 toxref = 4.23E-9 agidl = 7.698718012296599E-11
+ wagidl = 6.870229296090227E-17 bgidl = 1.52623582944205E9 wbgidl = -518.5486816927265
+ cgidl = 300 egidl = 0.1 noia = 1.5E42
+ noib = 0 noic = 0 em = 4.1E7
+ af = 1 ef = 1 kf = 0
+ lintnoi = -2E-7 tnoia = 2.5E7 tnoib = 0
+ ntnoi = 1 rnoia = 0.69 rnoib = 0.34
+ xpart = 0 cgso = {5.248925E-11/sw_func_tox_lv_ratio} cgdo = {5.248925E-11/sw_func_tox_lv_ratio}
+ cgbo = {0/sw_func_tox_lv_ratio} ckappas = 0.6 cf = 1.2E-11
+ clc = 1E-7 cle = 0.6 dlc = -3E-9
+ dwc = 0 vfbcv = -0.14469 noff = 3.9
+ voffcv = -0.10701 acde = 0.8 moin = 18.13
+ cgsl = {9.548271750000001E-12/sw_func_tox_lv_ratio} cgdl = {9.548271750000001E-12/sw_func_tox_lv_ratio} ijthsrev = 0.1
+ ijthsfwd = 0.1 xjbvs = 1 bvs = 12.69
+ jss = 2.1483E-5 jsws = 8.040000000000001E-10 cjs = {sw_psd_nw_cj}
+ mjs = 0.34629 mjsws = 0.29781 cjsws = {9.888891999999999E-11*sw_func_psd_nw_cj}
+ cjswgs = {2.39155046E-10*sw_func_psd_nw_cj} mjswgs = 0.9274 pbs = 0.6587
+ pbsws = 0.7418 pbswgs = 1.4338 xrcrg1 = 12
+ xrcrg2 = 1 rbpb = 50 rbpd = 50
+ rbps = 50 rbdb = 50 rbsb = 50
+ gbmin = 1E-12 tnom = 30 ute = 0.364939084399201
+ wute = -1.600709603142115E-6 kt1 = -0.39441525983983 wkt1 = -1.489861176348584E-7
+ kt1l = 0 kt2 = -0.05275360778419 wkt2 = 2.656694075999129E-10
+ ua1 = 3.27553940657852E-9 wua1 = -3.480000654845103E-15 ub1 = -1.345876590117556E-18
+ wub1 = 1.813335074212437E-24 uc1 = 1.61051151211626E-10 wuc1 = -1.506231605867368E-16
+ at = 1.29415688E5 wat = -0.117671287512834 prt = 0
+ njs = 1.3632 xtis = 5.2 tpb = 2.0386E-3
+ tpbsw = 1.246E-3 tpbswg = 0 tcj = 1.2407E-3
+ tcjsw = 3.7357E-4 tcjswg = 2E-12 tvoff = 0
+ tvfbsdoff = 0 saref = 3E-6 sbref = 3E-6
+ wlod = 0 ku0 = 4.5E-8 kvsat = 0.5
+ kvth0 = 3.29E-8 tku0 = 0 llodku0 = 0
+ wlodku0 = 1 llodvth = 0 wlodvth = 1
+ lku0 = 0 wku0 = 2.5E-7 pku0 = 0
+ lkvth0 = 0 wkvth0 = 2E-7 pkvth0 = 0
+ stk2 = 0 lodk2 = 1 steta0 = 0
+ lodeta0 = 1

.model pshort_model.26 pmos
+ level = 54 lmin = 4E-6 lmax = 8E-6 wmin = 1E-6
+ wmax = 3E-6 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 4.23E-9
+ toxm = 4.23E-9 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 9.999999999999999E22 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {7.3039E-9+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {-1.3994E-8-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = -5.722E-9 dwb = -1.7864E-8 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = -1.070590678651296 lvth0 = 7.236434194135481E-8
+ wvth0 = 5.332405039907553E-8 pvth0 = -9.73403684685344E-14 k1 = 0.319595437406316
+ lk1 = 5.584733025717702E-7 wk1 = 2.113469456509608E-7 pk1 = -8.849816241500118E-13
+ k2 = 0.058308404880749 lk2 = -2.015579481629036E-7 wk2 = -7.210020565219712E-8
+ pk2 = 2.948901581601409E-13 k3 = -15.845 k3b = 2
+ w0 = 0 lpe0 = 0 lpeb = 0
+ vbm = -3 dvtp0 = 0 dvtp1 = 0
+ dvt0 = 4.4955 dvt1 = 0.294 dvt2 = 0.015
+ dvt0w = -4.9772 dvt1w = 1.1472E6 dvt2w = -8.96E-3
+ vfbsdoff = 0 u0 = 0.015674420852953 lu0 = -1.192572203149783E-8
+ wu0 = -1.149947469000449E-8 pu0 = 2.937145862648324E-14 ua = 8.315481752881404E-10
+ lua = -3.414211394547378E-15 wua = -2.782795380006839E-15 pua = 7.959405580599845E-21
+ ub = 1.33704921227341E-19 lub = 2.185508852075004E-24 wub = 1.601206627797862E-24
+ pub = -5.227342987293764E-30 uc = -1.558841019870434E-10 luc = 2.237106289724087E-16
+ wuc = 1.307921533895637E-16 puc = -3.451437371283256E-22 ud = 0
+ up = 0 lp = 1 eu = 1.67
+ vsat = 8.185135232673584E4 lvsat = -0.235220972769428 wvsat = -0.013829074418523
+ pvsat = 1.322724154570256E-7 a0 = 1.045355568335618 la0 = 1.070606854900921E-7
+ wa0 = 2.411233684641524E-7 pa0 = -7.207799278397972E-13 ags = -0.092390242185578
+ lags = 1.784007885641172E-6 wags = 3.216187252773253E-7 pags = -1.330318646524736E-12
+ b0 = 0 b1 = 0 keta = 9.612565239788633E-3
+ lketa = -1.033745103942879E-7 wketa = 4.625743569724627E-10 pketa = 7.463765039419857E-14
+ a1 = 0 a2 = 0.8 rdsw = 547.88
+ rdswmin = 0 rdw = 0 rdwmin = 0
+ rsw = 0 rswmin = 0 prwb = -0.32348
+ prwg = 0.1376 wr = 1 voff = -0.248464494919859
+ lvoff = -3.324939584630798E-8 wvoff = -1.510061467262003E-8 pvoff = 1.224162945478934E-13
+ voffl = 0 minv = 0 nfactor = 2.122883907733277
+ lnfactor = -2.297426160838469E-6 wnfactor = -9.589219553653477E-7 pnfactor = 5.500664077226244E-12
+ eta0 = 0.08 etab = -0.07 dsub = 0.56
+ cit = 1E-5 cdsc = 1.3E-4 cdscb = 7.8E-4
+ cdscd = 0 pclm = -0.157542082732887 lpclm = 3.040636523860712E-6
+ wpclm = 1.20971853292584E-7 ppclm = -2.707342804998115E-12 pdiblc1 = 0.39
+ pdiblc2 = 2.051353797595502E-4 lpdiblc2 = -1.593344166247278E-9 wpdiblc2 = -1.090178070811516E-10
+ ppdiblc2 = 5.314502945718411E-15 pdiblcb = 0.07353922 wpdiblcb = -2.94178218782084E-7
+ drout = 0.56 pscbe1 = 6.715778682576205E8 lpscbe1 = 517.2828452842033
+ wpscbe1 = 126.51709511117947 ppscbe1 = -5.096094593973231E-4 pscbe2 = 9.344937673100734E-9
+ lpscbe2 = 6.864135332458846E-16 wpscbe2 = 2.665489798449702E-15 ppscbe2 = -1.078605020596392E-20
+ pvag = 0 delta = 0.01 fprout = 0
+ pdits = 0 pditsl = 0 pditsd = 0
+ lambda = 0 vtl = 0 lc = 5E-9
+ xn = 3 alpha0 = 3.148695103068001E-11 lalpha0 = -3.92835911380165E-17
+ walpha0 = -3.102699594741404E-17 palpha0 = 3.870974429539058E-23 alpha1 = -1.33069801511155E-12
+ lalpha1 = 1.068358332509587E-17 walpha1 = 1.311259444646403E-18 palpha1 = -1.052751967659953E-23
+ beta0 = 9.708507883125126 lbeta0 = -8.060528666919701E-5 wbeta0 = 1.999507805832999E-5
+ pbeta0 = 7.94278207625907E-11 aigbacc = 0.43 bigbacc = 0.054
+ cigbacc = 0.075 nigbacc = 1 aigbinv = 0.35
+ bigbinv = 0.03 cigbinv = 6E-3 eigbinv = 1.1
+ nigbinv = 3 aigc = 0.43 bigc = 0.054
+ cigc = 0.075 aigsd = 0.43 bigsd = 0.054
+ cigsd = 0.075 dlcig = 0 nigc = 1
+ poxedge = 1 pigcd = 1 ntox = 1
+ toxref = 4.23E-9 agidl = 2.861069588983125E-11 lagidl = 3.883658349057948E-16
+ wagidl = 1.056845273271772E-16 pagidl = -2.968929337056426E-22 bgidl = 2.056153730982706E9
+ lbgidl = -4.254174554553569E3 wbgidl = -1.040725648511257E3 pbgidl = 4.192030423495561E-3
+ cgidl = 300 egidl = 0.1 noia = 1.5E42
+ noib = 0 noic = 0 em = 4.1E7
+ af = 1 ef = 1 kf = 0
+ lintnoi = -2E-7 tnoia = 2.5E7 tnoib = 0
+ ntnoi = 1 rnoia = 0.69 rnoib = 0.34
+ xpart = 0 cgso = {5.248925E-11/sw_func_tox_lv_ratio} cgdo = {5.248925E-11/sw_func_tox_lv_ratio}
+ cgbo = {0/sw_func_tox_lv_ratio} ckappas = 0.6 cf = 1.2E-11
+ clc = 1E-7 cle = 0.6 dlc = -3E-9
+ dwc = 0 vfbcv = -0.14469 noff = 3.9
+ voffcv = -0.10701 acde = 0.8 moin = 18.13
+ cgsl = {9.548271750000001E-12/sw_func_tox_lv_ratio} cgdl = {9.548271750000001E-12/sw_func_tox_lv_ratio} ijthsrev = 0.1
+ ijthsfwd = 0.1 xjbvs = 1 bvs = 12.69
+ jss = 2.1483E-5 jsws = 8.040000000000001E-10 cjs = {sw_psd_nw_cj}
+ mjs = 0.34629 mjsws = 0.29781 cjsws = {9.888891999999999E-11*sw_func_psd_nw_cj}
+ cjswgs = {2.39155046E-10*sw_func_psd_nw_cj} mjswgs = 0.9274 pbs = 0.6587
+ pbsws = 0.7418 pbswgs = 1.4338 xrcrg1 = 12
+ xrcrg2 = 1 rbpb = 50 rbpd = 50
+ rbps = 50 rbdb = 50 rbsb = 50
+ gbmin = 1E-12 tnom = 30 ute = 0.931576961117328
+ lute = -4.548962074638601E-6 wute = -3.339395520765953E-6 pute = 1.395814968245316E-11
+ kt1 = -0.339727550906986 lkt1 = -4.390322710603627E-7 wkt1 = -2.865545212543623E-7
+ pkt1 = 1.104397493436534E-12 kt1l = 0 kt2 = -0.041841292291118
+ lkt2 = -8.760393783059053E-8 wkt2 = -3.603069283980048E-8 pkt2 = 2.913867605657834E-13
+ ua1 = 4.24753041995992E-9 lua1 = -7.803132191533705E-15 wua1 = -6.59666220600512E-15
+ pua1 = 2.5020521532774E-20 ub1 = -1.817318882535094E-18 lub1 = 3.784733066220485E-24
+ wub1 = 3.776085219719856E-24 pub1 = -1.575693461513182E-29 uc1 = 4.794595701344688E-10
+ luc1 = -2.556178966211554E-15 wuc1 = -3.768654827643817E-16 puc1 = 1.816270647534267E-21
+ at = 2.175299361574132E5 lat = -0.707380126836735 wat = -0.249417723927672
+ pat = 1.057658810581088E-6 prt = 0 njs = 1.3632
+ xtis = 5.2 tpb = 2.0386E-3 tpbsw = 1.246E-3
+ tpbswg = 0 tcj = 1.2407E-3 tcjsw = 3.7357E-4
+ tcjswg = 2E-12 tvoff = 0 tvfbsdoff = 0
+ saref = 3E-6 sbref = 3E-6 wlod = 0
+ ku0 = 4.5E-8 kvsat = 0.5 kvth0 = 3.29E-8
+ tku0 = 0 llodku0 = 0 wlodku0 = 1
+ llodvth = 0 wlodvth = 1 lku0 = 0
+ wku0 = 2.5E-7 pku0 = 0 lkvth0 = 0
+ wkvth0 = 2E-7 pkvth0 = 0 stk2 = 0
+ lodk2 = 1 steta0 = 0 lodeta0 = 1

.model pshort_model.27 pmos
+ level = 54 lmin = 2E-6 lmax = 4E-6 wmin = 1E-6
+ wmax = 3E-6 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 4.23E-9
+ toxm = 4.23E-9 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 9.999999999999999E22 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {7.3039E-9+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {-1.3994E-8-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = -5.722E-9 dwb = -1.7864E-8 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = -1.062589547191282 lvth0 = 4.013588043399419E-8
+ wvth0 = 3.596719676832147E-8 pvth0 = -2.74271703261006E-14 k1 = 0.376554545934803
+ lk1 = 3.290426969283286E-7 wk1 = 6.066643611828646E-8 pk1 = -2.780423399185139E-13
+ k2 = 0.038811895018855 lk2 = -1.230262403973134E-7 wk2 = -2.549804314202564E-8
+ pk2 = 1.071772067951203E-13 k3 = -15.845 k3b = 2
+ w0 = 0 lpe0 = 0 lpeb = 0
+ vbm = -3 dvtp0 = 0 dvtp1 = 0
+ dvt0 = 4.4955 dvt1 = 0.294 dvt2 = 0.015
+ dvt0w = -4.9772 dvt1w = 1.1472E6 dvt2w = -8.96E-3
+ vfbsdoff = 0 u0 = 0.015912534589053 lu0 = -1.288484130314656E-8
+ wu0 = -6.753727598515307E-9 pu0 = 1.025564629092992E-14 ua = 6.689537241546602E-10
+ lua = -2.759282896515133E-15 wua = -1.287505012169049E-15 pua = 1.936393922433641E-21
+ ub = 3.443428430135248E-19 lub = 1.337061830775318E-24 wub = 4.722331942566241E-25
+ pub = -6.798515446708609E-31 uc = -1.269527826910442E-10 luc = 1.071756220239558E-16
+ wuc = 6.179434897004269E-17 puc = -6.722140890014814E-23 ud = 0
+ up = 0 lp = 1 eu = 1.67
+ vsat = 3.667931015840721E4 lvsat = -0.053268528979907 wvsat = -4.705139586554242E-3
+ pvsat = 9.55213154410745E-8 a0 = 1.280594110078524 la0 = -8.404773377878359E-7
+ wa0 = -6.827138836937253E-8 pa0 = 5.254584399485593E-13 ags = 0.026539033954337
+ lags = 1.304962188500906E-6 wags = 2.110547138221196E-7 pags = -8.84968135151305E-13
+ b0 = 0 b1 = 0 keta = -1.756829069118203E-3
+ lketa = -5.757872655074284E-8 wketa = 1.293652676628547E-8 pketa = 2.439271977691468E-14
+ a1 = 0 a2 = 0.8 rdsw = 547.88
+ rdswmin = 0 rdw = 0 rdwmin = 0
+ rsw = 0 rswmin = 0 prwb = -0.32348
+ prwg = 0.1376 wr = 1 voff = -0.270487446847391
+ lvoff = 5.545879024236792E-8 wvoff = 3.212016373226919E-8 pvoff = -6.778843421765945E-14
+ voffl = 0 minv = 0 nfactor = 1.566782357526471
+ lnfactor = -5.7455789824058E-8 wnfactor = 6.951216060712303E-7 pnfactor = -1.161803539717556E-12
+ eta0 = 0.04028252430674 leta0 = 1.599815154827442E-7 weta0 = 1.185722421383489E-7
+ peta0 = -4.776075684663637E-13 etab = -0.035278433943364 letab = -1.398580514173367E-7
+ wetab = -1.036574924772655E-7 petab = 4.175311358085158E-13 dsub = 0.41012273323298
+ ldsub = 6.037038320103558E-7 wdsub = 4.474424231635809E-7 pdsub = -1.802292711193826E-12
+ cit = 1E-5 cdsc = 1.3E-4 cdscb = 7.8E-4
+ cdscd = 0 pclm = 0.749708856024025 lpclm = -6.137593704408655E-7
+ wpclm = -1.015335416706034E-6 ppclm = 1.869689242869078E-12 pdiblc1 = 0.39
+ pdiblc2 = -6.015393691001837E-4 lpdiblc2 = 1.655932042062744E-9 wpdiblc2 = 2.437690263504609E-9
+ ppdiblc2 = -4.943606602104185E-15 pdiblcb = 0.037724266543466 lpdiblcb = 1.442622027434792E-7
+ wpdiblcb = -2.58886443002652E-7 ppdiblcb = -1.42154849338243E-13 drout = 0.56
+ pscbe1 = 7.9999998E8 pscbe2 = 1.017347089412952E-8 lpscbe2 = -2.650908338659393E-15
+ wpscbe2 = -5.301553189921149E-16 ppscbe2 = 2.085969979350312E-21 pvag = 0
+ delta = 0.01 fprout = 0 pdits = 0
+ pditsl = 0 pditsd = 0 lambda = 0
+ vtl = 0 lc = 5E-9 xn = 3
+ alpha0 = -3.10384988888338E-11 lalpha0 = 2.125681708323861E-16 walpha0 = 2.753860245164431E-17
+ palpha0 = -1.971917832688357E-22 alpha1 = -1.486981758121058E-10 lalpha1 = 6.042780154816553E-16
+ walpha1 = 1.465289440676121E-16 palpha1 = -5.954626107256897E-22 beta0 = -29.114678942622973
+ lbeta0 = 7.577404398667438E-5 wbeta0 = 8.522905155362852E-5 pbeta0 = -1.833338416687898E-10
+ aigbacc = 0.43 bigbacc = 0.054 cigbacc = 0.075
+ nigbacc = 1 aigbinv = 0.35 bigbinv = 0.03
+ cigbinv = 6E-3 eigbinv = 1.1 nigbinv = 3
+ aigc = 0.43 bigc = 0.054 cigc = 0.075
+ aigsd = 0.43 bigsd = 0.054 cigsd = 0.075
+ dlcig = 0 nigc = 1 poxedge = 1
+ pigcd = 1 ntox = 1 toxref = 4.23E-9
+ agidl = 1.353662280421619E-10 lagidl = -4.164416753740723E-17 wagidl = -6.90401414974663E-17
+ pagidl = 4.068959356239955E-22 bgidl = 1E9 cgidl = 300
+ egidl = 0.1 noia = 1.5E42 noib = 0
+ noic = 0 em = 4.1E7 af = 1
+ ef = 1 kf = 0 lintnoi = -2E-7
+ tnoia = 2.5E7 tnoib = 0 ntnoi = 1
+ rnoia = 0.69 rnoib = 0.34 xpart = 0
+ cgso = {5.248925E-11/sw_func_tox_lv_ratio} cgdo = {5.248925E-11/sw_func_tox_lv_ratio} cgbo = {0/sw_func_tox_lv_ratio}
+ ckappas = 0.6 cf = 1.2E-11 clc = 1E-7
+ cle = 0.6 dlc = -3E-9 dwc = 0
+ vfbcv = -0.14469 noff = 3.9 voffcv = -0.10701
+ acde = 0.8 moin = 18.13 cgsl = {9.548271750000001E-12/sw_func_tox_lv_ratio}
+ cgdl = {9.548271750000001E-12/sw_func_tox_lv_ratio} ijthsrev = 0.1 ijthsfwd = 0.1
+ xjbvs = 1 bvs = 12.69 jss = 2.1483E-5
+ jsws = 8.040000000000001E-10 cjs = {sw_psd_nw_cj} mjs = 0.34629
+ mjsws = 0.29781 cjsws = {9.888891999999999E-11*sw_func_psd_nw_cj} cjswgs = {2.39155046E-10*sw_func_psd_nw_cj}
+ mjswgs = 0.9274 pbs = 0.6587 pbsws = 0.7418
+ pbswgs = 1.4338 xrcrg1 = 12 xrcrg2 = 1
+ rbpb = 50 rbpd = 50 rbps = 50
+ rbdb = 50 rbsb = 50 gbmin = 1E-12
+ tnom = 30 ute = 0.73942528501565 lute = -3.774977429121153E-6
+ wute = 2.677356397033453E-8 pute = 3.99261003164412E-13 kt1 = -0.420624909816988
+ lkt1 = -1.131786801391806E-7 wkt1 = -3.037913732348676E-8 pkt1 = 7.252612106757463E-14
+ kt1l = 0 kt2 = -0.065750969778062 lkt2 = 8.703956170688232E-9
+ wkt2 = 5.721076262101811E-8 pkt2 = -8.418870313292837E-14 ua1 = 4.842536580090784E-9
+ lua1 = -1.019980986446691E-14 wua1 = -8.090250067559783E-16 pua1 = 1.707988345844845E-21
+ ub1 = -2.325048766884653E-18 lub1 = 5.829862947621896E-24 wub1 = -4.703289977534112E-25
+ pub1 = 1.347570895879896E-30 uc1 = -2.968448437955069E-10 luc1 = 5.707658974454206E-16
+ wuc1 = 7.192729550517714E-17 puc1 = 8.538722177823065E-24 at = 4.693175886721143E4
+ lat = -0.02021271588993 wat = 0.055984841331432 pat = -1.724990574518011E-7
+ prt = 0 njs = 1.3632 xtis = 5.2
+ tpb = 2.0386E-3 tpbsw = 1.246E-3 tpbswg = 0
+ tcj = 1.2407E-3 tcjsw = 3.7357E-4 tcjswg = 2E-12
+ tvoff = 0 tvfbsdoff = 0 saref = 3E-6
+ sbref = 3E-6 wlod = 0 ku0 = 4.5E-8
+ kvsat = 0.5 kvth0 = 3.29E-8 tku0 = 0
+ llodku0 = 0 wlodku0 = 1 llodvth = 0
+ wlodvth = 1 lku0 = 0 wku0 = 2.5E-7
+ pku0 = 0 lkvth0 = 0 wkvth0 = 2E-7
+ pkvth0 = 0 stk2 = 0 lodk2 = 1
+ steta0 = 0 lodeta0 = 1

.model pshort_model.28 pmos
+ level = 54 lmin = 1E-6 lmax = 2E-6 wmin = 1E-6
+ wmax = 3E-6 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 4.23E-9
+ toxm = 4.23E-9 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 9.999999999999999E22 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {7.3039E-9+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {-1.3994E-8-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = -5.722E-9 dwb = -1.7864E-8 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = -1.070583647158006 lvth0 = 5.634781923731091E-8
+ wvth0 = 4.04840108665631E-8 pvth0 = -3.658721511556546E-14 k1 = 0.584693988804693
+ lk1 = -9.30615955384937E-8 wk1 = -1.139299673479209E-7 pk1 = 7.603707115411307E-14
+ k2 = -0.042980437511446 lk2 = 4.284762846614701E-8 wk2 = 4.656228443579386E-8
+ pk2 = -3.896027280876672E-14 k3 = -15.845 k3b = 2
+ w0 = 0 lpe0 = 0 lpeb = 0
+ vbm = -3 dvtp0 = 0 dvtp1 = 0
+ dvt0 = 4.4955 dvt1 = 0.294 dvt2 = 0.015
+ dvt0w = -4.9772 dvt1w = 1.1472E6 dvt2w = -8.96E-3
+ vfbsdoff = 0 u0 = 0.013569861178814 lu0 = -8.13392773926149E-9
+ wu0 = -6.471148461236285E-9 pu0 = 9.68257919147771E-15 ua = 2.914734354092558E-10
+ lua = -1.993757400702918E-15 wua = -1.567223836744917E-15 pua = 2.503660342047606E-21
+ ub = 4.222846579752419E-19 lub = 1.178996765334735E-24 wub = 8.879995402590949E-25
+ pub = -1.523020705167719E-30 uc = -1.287555144549242E-10 luc = 1.108315404083232E-16
+ wuc = 8.619486387220365E-17 puc = -1.167053603155518E-22 ud = 0
+ up = 0 lp = 1 eu = 1.67
+ vsat = -8.519367640077221E4 lvsat = 0.193888425286271 wvsat = 0.161552382679402
+ pvsat = -2.416469446240184E-7 a0 = 0.422167560128885 la0 = 9.004014043914338E-7
+ wa0 = 1.143223087814755E-6 pa0 = -1.931437819819138E-12 ags = 1.001545272866255
+ lags = -6.723387639375953E-7 wags = -1.355994578433244E-6 pags = 2.292989024951066E-12
+ b0 = 0 b1 = 0 keta = -0.068167309744583
+ lketa = 7.710093133333258E-8 wketa = 9.588254661323742E-8 pketa = -1.438208131204657E-13
+ a1 = 0 a2 = 0.8 rdsw = 547.88
+ rdswmin = 0 rdw = 0 rdwmin = 0
+ rsw = 0 rswmin = 0 prwb = -0.32348
+ prwg = 0.1376 wr = 1 voff = -0.229915733566203
+ lvoff = -2.682015743132242E-8 wvoff = -1.649147786522788E-8 pvoff = 3.079539160236544E-14
+ voffl = 0 minv = 0 nfactor = 1.971454968599019
+ lnfactor = -8.781269890078523E-7 wnfactor = -4.640419309881576E-7 pnfactor = 1.188966203476438E-12
+ eta0 = -0.469699256776667 leta0 = 1.194218447738521E-6 weta0 = 3.827994572004839E-7
+ peta0 = -1.013457189885793E-12 etab = 34.730508313192715 letab = -7.064445638516834E-5
+ wetab = -3.421708037911301E-5 petab = 6.959914338883118E-11 dsub = 1.32009663706808
+ ldsub = -1.241712325280382E-6 wdsub = -1.348502364481197E-6 pdsub = 1.839861766812332E-12
+ cit = 1E-5 cdsc = 1.3E-4 cdscb = 7.8E-4
+ cdscd = 0 pclm = 0.132614860746103 lpclm = 6.376998468548167E-7
+ wpclm = 1.971269652867263E-7 ppclm = -5.891699182636558E-13 pdiblc1 = 0.407396735930792
+ lpdiblc1 = -3.528037170681464E-8 wpdiblc1 = -9.281271471358518E-9 ppdiblc1 = 1.882230716865742E-14
+ pdiblc2 = -1.149118408660619E-4 lpdiblc2 = 6.690572543342833E-10 wpdiblc2 = 3.250925546770588E-10
+ ppdiblc2 = -6.592837997744191E-16 pdiblcb = 0.209296854858191 lpdiblcb = -2.036849474877231E-7
+ wpdiblcb = -6.305470046405131E-7 ppdiblcb = 6.115683097365995E-13 drout = 0.431913827537372
+ ldrout = 2.597572207201402E-7 wdrout = -2.295939101561477E-7 pdrout = 4.656136946697457E-13
+ pscbe1 = 8E8 pscbe2 = 1.093508405381235E-8 lpscbe2 = -4.19545068713827E-15
+ wpscbe2 = -5.653620751791414E-16 ppscbe2 = 2.157368858416528E-21 pvag = 0
+ delta = 0.01 fprout = 0 pdits = 0
+ pditsl = 0 pditsd = 0 lambda = 0
+ vtl = 0 lc = 5E-9 xn = 3
+ alpha0 = 4.68236675478178E-11 lalpha0 = 5.46646316448539E-17 walpha0 = -1.413438279601305E-16
+ palpha0 = 1.452997590170786E-22 alpha1 = 1.999210993128143E-10 lalpha1 = -1.027176910403814E-16
+ walpha1 = -2.983036705039013E-16 palpha1 = 3.066525936339644E-22 beta0 = 7.616416095732391
+ lbeta0 = 1.283824022030168E-6 wbeta0 = -1.052655092956784E-5 pbeta0 = 1.085737109990262E-11
+ aigbacc = 0.43 bigbacc = 0.054 cigbacc = 0.075
+ nigbacc = 1 aigbinv = 0.35 bigbinv = 0.03
+ cigbinv = 6E-3 eigbinv = 1.1 nigbinv = 3
+ aigc = 0.43 bigc = 0.054 cigc = 0.075
+ aigsd = 0.43 bigsd = 0.054 cigsd = 0.075
+ dlcig = 0 nigc = 1 poxedge = 1
+ pigcd = 1 ntox = 1 toxref = 4.23E-9
+ agidl = 1.300781185373606E-10 lagidl = -3.091994491898421E-17 wagidl = 2.668833571488318E-16
+ pagidl = -2.743528885487133E-22 bgidl = 6.955255896436541E8 lbgidl = 617.4704505097452
+ wbgidl = 300.0267090647425 pbgidl = -6.084505656627889E-4 cgidl = 300
+ egidl = 0.1 noia = 1.5E42 noib = 0
+ noic = 0 em = 4.1E7 af = 1
+ ef = 1 kf = 0 lintnoi = -2E-7
+ tnoia = 2.5E7 tnoib = 0 ntnoi = 1
+ rnoia = 0.69 rnoib = 0.34 xpart = 0
+ cgso = {5.248925E-11/sw_func_tox_lv_ratio} cgdo = {5.248925E-11/sw_func_tox_lv_ratio} cgbo = {0/sw_func_tox_lv_ratio}
+ ckappas = 0.6 cf = 1.2E-11 clc = 1E-7
+ cle = 0.6 dlc = -3E-9 dwc = 0
+ vfbcv = -0.14469 noff = 3.9 voffcv = -0.10701
+ acde = 0.8 moin = 18.13 cgsl = {9.548271750000001E-12/sw_func_tox_lv_ratio}
+ cgdl = {9.548271750000001E-12/sw_func_tox_lv_ratio} ijthsrev = 0.1 ijthsfwd = 0.1
+ xjbvs = 1 bvs = 12.69 jss = 2.1483E-5
+ jsws = 8.040000000000001E-10 cjs = {sw_psd_nw_cj} mjs = 0.34629
+ mjsws = 0.29781 cjsws = {9.888891999999999E-11*sw_func_psd_nw_cj} cjswgs = {2.39155046E-10*sw_func_psd_nw_cj}
+ mjswgs = 0.9274 pbs = 0.6587 pbsws = 0.7418
+ pbswgs = 1.4338 xrcrg1 = 12 xrcrg2 = 1
+ rbpb = 50 rbpd = 50 rbps = 50
+ rbdb = 50 rbsb = 50 gbmin = 1E-12
+ tnom = 30 ute = -2.255587171094037 lute = 2.298871891719819E-6
+ wute = 1.642914629133077E-6 pute = -2.878253683292849E-12 kt1 = -0.536572938317938
+ lkt1 = 1.219625302844033E-7 wkt1 = 1.080775230828379E-7 pkt1 = -2.082623247565268E-13
+ kt1l = 0 kt2 = -0.079967295607865 lkt2 = 3.753449435761798E-8
+ wkt2 = 5.25196157051104E-8 pkt2 = -7.467511348123053E-14 ua1 = -8.879427949752057E-10
+ lua1 = 1.421533542414418E-15 wua1 = 8.121843413064413E-16 pua1 = -1.579804757513565E-21
+ ub1 = 5.713159946608073E-19 lub1 = -4.393003241515891E-26 wub1 = 4.430427686762031E-25
+ pub1 = -5.047360859781646E-31 uc1 = -1.521523209212733E-10 luc1 = 2.773311973667494E-16
+ wuc1 = 2.255085773013926E-16 puc1 = -3.029222743295203E-22 at = -1.283494791995439E4
+ lat = 0.100993448273961 wat = 4.306496088416198E-3 pat = -6.769599343910778E-8
+ prt = 0 njs = 1.3632 xtis = 5.2
+ tpb = 2.0386E-3 tpbsw = 1.246E-3 tpbswg = 0
+ tcj = 1.2407E-3 tcjsw = 3.7357E-4 tcjswg = 2E-12
+ tvoff = 0 tvfbsdoff = 0 saref = 3E-6
+ sbref = 3E-6 wlod = 0 ku0 = 4.5E-8
+ kvsat = 0.5 kvth0 = 3.29E-8 tku0 = 0
+ llodku0 = 0 wlodku0 = 1 llodvth = 0
+ wlodvth = 1 lku0 = 0 wku0 = 2.5E-7
+ pku0 = 0 lkvth0 = 0 wkvth0 = 2E-7
+ pkvth0 = 0 stk2 = 0 lodk2 = 1
+ steta0 = 0 lodeta0 = 1

.model pshort_model.29 pmos
+ level = 54 lmin = 5E-7 lmax = 1E-6 wmin = 1E-6
+ wmax = 3E-6 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 4.23E-9
+ toxm = 4.23E-9 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 9.999999999999999E22 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {7.3039E-9+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {-1.3994E-8-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = -5.722E-9 dwb = -1.7864E-8 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = -1.037206619589629 lvth0 = 2.203663542135025E-8
+ wvth0 = -6.799919121476631E-9 pvth0 = 1.202009750497953E-14 k1 = 0.570478311334409
+ lk1 = -7.844804968717182E-8 wk1 = -1.729151313343002E-7 pk1 = 1.366731119101431E-13
+ k2 = -0.032483973546996 lk2 = 3.205738946826014E-8 wk2 = 5.39584854093795E-8
+ pk2 = -4.656347865520108E-14 k3 = -15.845 k3b = 2
+ w0 = 0 lpe0 = 0 lpeb = 0
+ vbm = -3 dvtp0 = 0 dvtp1 = 0
+ dvt0 = 4.4955 dvt1 = 0.294 dvt2 = 0.015
+ dvt0w = -4.9772 dvt1w = 1.1472E6 dvt2w = -8.96E-3
+ vfbsdoff = 0 u0 = 4.132218653956039E-3 lu0 = 1.567855524581807E-9
+ wu0 = 6.172387042884386E-9 pu0 = -3.31482358433229E-15 ua = -2.071001846484218E-9
+ lua = 4.348388393801906E-16 wua = 1.670041410082155E-15 pua = -8.242094845076614E-22
+ ub = 1.840578805828502E-18 lub = -2.789925991286426E-25 wub = -1.121231636192164E-24
+ pub = 5.424448334500571E-31 uc = -4.311489715324689E-11 luc = 2.279401350960657E-17
+ wuc = -3.34564346762489E-17 puc = 6.294738776674884E-24 ud = 0
+ up = 0 lp = 1 eu = 1.67
+ vsat = 1.177275056360264E5 lvsat = -0.014712114793374 wvsat = -0.151256346740628
+ pvsat = 7.991667551502013E-8 a0 = 1.675147541233958 la0 = -3.876469804248083E-7
+ wa0 = -1.714666393775812E-6 pa0 = 1.006438272582186E-12 ags = -0.182888202294138
+ lags = 5.452446353255858E-7 wags = 1.316446917063464E-6 pags = -4.542487631216037E-13
+ b0 = 0 b1 = 0 keta = 0.016237083599563
+ lketa = -9.665772171730056E-9 wketa = -5.795371406290034E-8 pketa = 1.432101681947578E-14
+ a1 = 0 a2 = 0.735070884838401 la2 = 6.674635123674226E-8
+ wa2 = 6.398064363314183E-8 pa2 = -6.577133388714618E-14 rdsw = 547.88
+ rdswmin = 0 rdw = 0 rdwmin = 0
+ rsw = 0 rswmin = 0 prwb = -0.32348
+ prwg = 0.1376 wr = 1 voff = -0.249376219748871
+ lvoff = -6.815011161374093E-9 wvoff = 7.509121956665707E-9 pvoff = 6.123062992656693E-15
+ voffl = 0 minv = 0 nfactor = 0.88972097903658
+ lnfactor = 2.3388257145446E-7 wnfactor = 8.3516165461627E-7 pnfactor = -1.465994920818866E-13
+ eta0 = 0.905318256326376 leta0 = -2.192830555212506E-7 weta0 = -1.239887882954364E-6
+ peta0 = 6.546459235453084E-13 etab = -69.88309008149675 letab = 3.689706740139167E-5
+ wetab = 6.884807678264845E-5 petab = -3.635060139157366E-11 dsub = -0.06024441375882
+ ldsub = 1.772617108770616E-7 wdsub = 8.636023326827938E-7 pdsub = -4.341553166158842E-13
+ cit = 1E-5 cdsc = 1.3E-4 cdscb = 7.8E-4
+ cdscd = 0 pclm = 0.892106295025021 lpclm = -1.430482336866988E-7
+ wpclm = -7.783078756765857E-7 ppclm = 4.135653930285371E-13 pdiblc1 = 0.549646572599227
+ lpdiblc1 = -1.815114968039257E-7 wpdiblc1 = 7.133441101795747E-8 ppdiblc1 = -6.404964704216953E-14
+ pdiblc2 = 4.528330516008606E-4 lpdiblc2 = 8.542231781699661E-11 wpdiblc2 = -5.644133926565035E-10
+ ppdiblc2 = 2.551176400131148E-16 pdiblcb = 0.364589066867197 lpdiblcb = -3.633234779264375E-7
+ wpdiblcb = -3.838980276962143E-7 ppdiblcb = 3.580161212255837E-13 drout = 0.351542904925256
+ ldrout = 3.423775647143237E-7 wdrout = 4.591878203122953E-7 pdrout = -2.424456588710482E-13
+ pscbe1 = 8E8 pscbe2 = 4.24306980430433E-9 lpscbe2 = 2.683859657184982E-15
+ wpscbe2 = 3.161837807944958E-15 ppscbe2 = -1.674147895036448E-21 pvag = 0
+ delta = 0.01 fprout = 0 pdits = 0
+ pditsl = 0 pditsd = 0 lambda = 0
+ vtl = 0 lc = 5E-9 xn = 3
+ alpha0 = 1E-10 alpha1 = 1E-10 beta0 = 8.130897551755378
+ lbeta0 = 7.549432590160084E-7 wbeta0 = 6.227142997885776E-7 pbeta0 = -6.039397646930265E-13
+ aigbacc = 0.43 bigbacc = 0.054 cigbacc = 0.075
+ nigbacc = 1 aigbinv = 0.35 bigbinv = 0.03
+ cigbinv = 6E-3 eigbinv = 1.1 nigbinv = 3
+ aigc = 0.43 bigc = 0.054 cigc = 0.075
+ aigsd = 0.43 bigsd = 0.054 cigsd = 0.075
+ dlcig = 0 nigc = 1 poxedge = 1
+ pigcd = 1 ntox = 1 toxref = 4.23E-9
+ agidl = 7.528645472124368E-11 lagidl = 2.540522798401818E-17 wagidl = -2.653003610458662E-16
+ pagidl = 2.727255875508179E-22 bgidl = 1.608948820712692E9 lbgidl = -321.51766995045267
+ wbgidl = -600.053418129485 pbgidl = 3.168210041313504E-4 cgidl = 300
+ egidl = 0.1 noia = 1.5E42 noib = 0
+ noic = 0 em = 4.1E7 af = 1
+ ef = 1 kf = 0 lintnoi = -2E-7
+ tnoia = 2.5E7 tnoib = 0 ntnoi = 1
+ rnoia = 0.69 rnoib = 0.34 xpart = 0
+ cgso = {5.248925E-11/sw_func_tox_lv_ratio} cgdo = {5.248925E-11/sw_func_tox_lv_ratio} cgbo = {0/sw_func_tox_lv_ratio}
+ ckappas = 0.6 cf = 1.2E-11 clc = 1E-7
+ cle = 0.6 dlc = -3E-9 dwc = 0
+ vfbcv = -0.14469 noff = 3.9 voffcv = -0.10701
+ acde = 0.8 moin = 18.13 cgsl = {9.548271750000001E-12/sw_func_tox_lv_ratio}
+ cgdl = {9.548271750000001E-12/sw_func_tox_lv_ratio} ijthsrev = 0.1 ijthsfwd = 0.1
+ xjbvs = 1 bvs = 12.69 jss = 2.1483E-5
+ jsws = 8.040000000000001E-10 cjs = {sw_psd_nw_cj} mjs = 0.34629
+ mjsws = 0.29781 cjsws = {9.888891999999999E-11*sw_func_psd_nw_cj} cjswgs = {2.39155046E-10*sw_func_psd_nw_cj}
+ mjswgs = 0.9274 pbs = 0.6587 pbsws = 0.7418
+ pbswgs = 1.4338 xrcrg1 = 12 xrcrg2 = 1
+ rbpb = 50 rbpd = 50 rbps = 50
+ rbdb = 50 rbsb = 50 gbmin = 1E-12
+ tnom = 30 ute = 0.335781545423211 lute = -3.650240524353136E-7
+ wute = -2.498312697460492E-6 pute = 1.378878313717421E-12 kt1 = -0.322334465902354
+ lkt1 = -9.82720484971478E-8 wkt1 = -1.943198559152932E-7 pkt1 = 1.025985520850038E-13
+ kt1l = 0 kt2 = -0.031064648351439 lkt2 = -1.273684019022031E-8
+ wkt2 = -4.137115754353098E-8 pkt2 = 2.184347472909383E-14 ua1 = 4.301335980268917E-10
+ lua1 = 6.656682732497756E-17 wua1 = -1.489778001725278E-15 pua1 = 7.865849075749257E-22
+ ub1 = 7.158246909607063E-19 lub1 = -1.924832381070996E-25 wub1 = -3.069520994055133E-25
+ pub1 = 2.662496384714229E-31 uc1 = 2.161595382550631E-10 luc1 = -1.012889741242142E-16
+ wuc1 = -1.422043259332327E-16 puc1 = 7.508217764083567E-23 at = 9.296300050203098E4
+ lat = -7.765573128458741E-3 wat = -0.112745290115544 pat = 5.263183815712845E-8
+ prt = 0 njs = 1.3632 xtis = 5.2
+ tpb = 2.0386E-3 tpbsw = 1.246E-3 tpbswg = 0
+ tcj = 1.2407E-3 tcjsw = 3.7357E-4 tcjswg = 2E-12
+ tvoff = 0 tvfbsdoff = 0 saref = 2.75E-6
+ sbref = 2.74E-6 wlod = 0 ku0 = 4.5E-8
+ kvsat = 0.5 kvth0 = 3.29E-8 tku0 = 0
+ llodku0 = 0 wlodku0 = 1 llodvth = 0
+ wlodvth = 1 lku0 = 0 wku0 = 2.5E-7
+ pku0 = 0 lkvth0 = 0 wkvth0 = 2E-7
+ pkvth0 = 0 stk2 = 0 lodk2 = 1
+ steta0 = 0 lodeta0 = 1

.model pshort_model.30 pmos
+ level = 54 lmin = 2.5E-7 lmax = 5E-7 wmin = 1E-6
+ wmax = 3E-6 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 4.23E-9
+ toxm = 4.23E-9 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 9.999999999999999E22 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {7.3039E-9+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {-1.3994E-8-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = -5.722E-9 dwb = -1.7864E-8 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = -1.004292618966362 lvth0 = 4.658438060272544E-9
+ wvth0 = 1.466828093097363E-8 pvth0 = 6.851454956864196E-16 k1 = -0.070397138826865
+ lk1 = 2.599264974925788E-7 wk1 = 4.931070937694629E-7 pk1 = -2.149786306779425E-13
+ k2 = 0.197642966135991 lk2 = -8.944687316108119E-8 wk2 = -1.846571049983218E-7
+ pk2 = 7.942268969298027E-14 k3 = -15.845 k3b = 2
+ w0 = 0 lpe0 = 0 lpeb = 0
+ vbm = -3 dvtp0 = 0 dvtp1 = 0
+ dvt0 = 4.4955 dvt1 = 0.294 dvt2 = 0.015
+ dvt0w = -4.9772 dvt1w = 1.1472E6 dvt2w = -8.96E-3
+ vfbsdoff = 0 u0 = 0.010538038403274 lu0 = -1.814340433220872E-9
+ wu0 = -1.259685690175206E-9 pu0 = 6.092216338503777E-16 ua = -2.543721792798865E-10
+ lua = -5.243198253476902E-16 wua = -3.651118545274771E-16 pua = 2.503270173670489E-22
+ ub = 6.184739807392808E-19 lub = 3.662640832605652E-25 wub = 2.32631393391777E-25
+ pub = -1.723785998139085E-31 uc = 1.082825524715168E-11 luc = -5.687323639975068E-18
+ wuc = -5.60925292486559E-17 puc = 1.824632507777091E-23 ud = 0
+ up = 0 lp = 1 eu = 1.67
+ vsat = 6.337643704419064E4 lvsat = 0.013984597210292 wvsat = -0.068595297839392
+ pvsat = 3.627263362775436E-8 a0 = 1.600747695555484 la0 = -3.48364754704722E-7
+ wa0 = -1.045263927245778E-7 pa0 = 1.563036737071474E-13 ags = 0.524354077808333
+ lags = 1.718291983388428E-7 wags = 1.752919761635912E-6 pags = -6.847011873817216E-13
+ b0 = 0 b1 = 0 keta = 0.118112293952102
+ lketa = -6.345466073534625E-8 wketa = -1.748817941936045E-7 pketa = 7.6057639991526E-14
+ a1 = 0 a2 = 0.77849879888746 la2 = 4.381693375380741E-8
+ wa2 = 3.239059787384056E-7 pa2 = -2.030087917187042E-13 rdsw = 547.88
+ rdswmin = 0 rdw = 0 rdwmin = 0
+ rsw = 0 rswmin = 0 prwb = -0.32348
+ prwg = 0.1376 wr = 1 voff = -0.220161396589751
+ lvoff = -2.224008721151149E-8 wvoff = 2.416298647595361E-8 pvoff = -2.669977627153084E-15
+ voffl = 0 minv = 0 nfactor = 0.815837240464689
+ lnfactor = 2.728922988155554E-7 wnfactor = 1.095243650171679E-6 pnfactor = -2.839196647511957E-13
+ eta0 = 0.817165172536417 leta0 = -1.727392851171578E-7 weta0 = -3.223860091290397E-7
+ peta0 = 1.702159441880234E-13 etab = -1.413508598212978E-3 letab = 3.807510201293091E-10
+ wetab = 1.448335267613062E-9 petab = -4.077308979529652E-16 dsub = 0.092847434604701
+ ldsub = 9.643105204330291E-8 wdsub = -1.190166744226618E-7 pdsub = 8.465572770771101E-14
+ cit = 1E-5 cdsc = 1.3E-4 cdscb = 7.8E-4
+ cdscd = 0 pclm = 0.251666451194038 lpclm = 1.950963185779337E-7
+ wpclm = 3.57116938528523E-7 ppclm = -1.859252837739896E-13 pdiblc1 = 0.045206262141436
+ lpdiblc1 = 8.482693383406247E-8 wpdiblc1 = -2.27822672428193E-7 ppdiblc1 = 9.39017031323966E-14
+ pdiblc2 = -5.533424091727651E-3 lpdiblc2 = 3.24609425440873E-9 wpdiblc2 = -5.566546354774411E-9
+ ppdiblc2 = 2.896183818415825E-15 pdiblcb = -0.599496649794652 lpdiblcb = 1.457022114424186E-7
+ wpdiblcb = 7.852462831486615E-7 ppdiblcb = -2.592780451687805E-13 drout = 1.375949172796848
+ ldrout = -1.984966518466621E-7 wdrout = 2.522563076572365E-7 pdrout = -1.33188303367329E-13
+ pscbe1 = 8E8 pscbe2 = 9.42793283167796E-9 lpscbe2 = -5.368580291196584E-17
+ wpscbe2 = 8.602245812576025E-18 ppscbe2 = -9.277357057296353E-24 pvag = 0
+ delta = 0.01 fprout = 0 pdits = 0
+ pditsl = 0 pditsd = 0 lambda = 0
+ vtl = 0 lc = 5E-9 xn = 3
+ alpha0 = 1E-10 alpha1 = 1E-10 beta0 = 10.473324426420923
+ lbeta0 = -4.818300216849029E-7 wbeta0 = -1.706669125818473E-6 pbeta0 = 6.259467314263892E-13
+ aigbacc = 0.43 bigbacc = 0.054 cigbacc = 0.075
+ nigbacc = 1 aigbinv = 0.35 bigbinv = 0.03
+ cigbinv = 6E-3 eigbinv = 1.1 nigbinv = 3
+ aigc = 0.43 bigc = 0.054 cigc = 0.075
+ aigsd = 0.43 bigsd = 0.054 cigsd = 0.075
+ dlcig = 0 nigc = 1 poxedge = 1
+ pigcd = 1 ntox = 1 toxref = 4.23E-9
+ agidl = -3.938494523778692E-9 lagidl = 2.144633419260243E-15 wagidl = 4.558806795070038E-15
+ pagidl = -2.274345101592506E-21 bgidl = 1.151951147073894E9 lbgidl = -80.22838224125098
+ wbgidl = -453.6337692554552 pbgidl = 2.395131865616492E-4 cgidl = 697.0613816756013
+ lcgidl = -2.096436447881373E-4 wcgidl = -3.912611884243604E-4 pcgidl = 2.065812123538012E-10
+ egidl = -2.001119726620334 legidl = 1.109366002218817E-6 wegidl = 2.07042698987781E-6
+ pegidl = -1.093160605531605E-12 noia = 1.5E42 noib = 0
+ noic = 0 em = 4.1E7 af = 1
+ ef = 1 kf = 0 lintnoi = -2E-7
+ tnoia = 2.5E7 tnoib = 0 ntnoi = 1
+ rnoia = 0.69 rnoib = 0.34 xpart = 0
+ cgso = {5.248925E-11/sw_func_tox_lv_ratio} cgdo = {5.248925E-11/sw_func_tox_lv_ratio} cgbo = {0/sw_func_tox_lv_ratio}
+ ckappas = 0.6 cf = 1.2E-11 clc = 1E-7
+ cle = 0.6 dlc = -3E-9 dwc = 0
+ vfbcv = -0.14469 noff = 3.9 voffcv = -0.10701
+ acde = 0.8 moin = 18.13 cgsl = {9.548271750000001E-12/sw_func_tox_lv_ratio}
+ cgdl = {9.548271750000001E-12/sw_func_tox_lv_ratio} ijthsrev = 0.1 ijthsfwd = 0.1
+ xjbvs = 1 bvs = 12.69 jss = 2.1483E-5
+ jsws = 8.040000000000001E-10 cjs = {sw_psd_nw_cj} mjs = 0.34629
+ mjsws = 0.29781 cjsws = {9.888891999999999E-11*sw_func_psd_nw_cj} cjswgs = {2.39155046E-10*sw_func_psd_nw_cj}
+ mjswgs = 0.9274 pbs = 0.6587 pbsws = 0.7418
+ pbswgs = 1.4338 xrcrg1 = 12 xrcrg2 = 1
+ rbpb = 50 rbpd = 50 rbps = 50
+ rbdb = 50 rbsb = 50 gbmin = 1E-12
+ tnom = 30 ute = -0.354500766427809 lute = -5.632751657175898E-10
+ wute = 5.154892435146603E-8 pute = 3.258197574016943E-14 kt1 = -0.467730935407027
+ lkt1 = -2.150445735631459E-8 wkt1 = -3.617859369566812E-8 pkt1 = 1.910186332818842E-14
+ kt1l = 0 kt2 = -0.025186402318738 lkt2 = -1.584048355653408E-8
+ wkt2 = -7.075760942414067E-8 pkt2 = 3.735916868463318E-14 ua1 = 1.06005742850985E-9
+ lua1 = -2.660253960840589E-16 wua1 = -3.281097505103061E-16 pua1 = 1.732380109524355E-22
+ ub1 = 3.305565442537945E-19 lub1 = 1.093372013638933E-26 wub1 = 3.41004012045752E-25
+ pub1 = -7.586341290150767E-32 uc1 = 5.067960087402845E-11 luc1 = -1.391755294627653E-17
+ wuc1 = 4.597559985466674E-20 puc1 = -2.427456501606578E-26 at = 1.084380419738865E5
+ lat = -0.015936209325101 wat = -0.044508430680046 pat = 1.660359521749901E-8
+ prt = 0 njs = 1.3632 xtis = 5.2
+ tpb = 2.0386E-3 tpbsw = 1.246E-3 tpbswg = 0
+ tcj = 1.2407E-3 tcjsw = 3.7357E-4 tcjswg = 2E-12
+ tvoff = 0 tvfbsdoff = 0 saref = 1.75E-6
+ sbref = 1.74E-6 wlod = 0 ku0 = 4.5E-8
+ kvsat = 0.5 kvth0 = 3.29E-8 tku0 = 0
+ llodku0 = 0 wlodku0 = 1 llodvth = 0
+ wlodvth = 1 lku0 = 0 wku0 = 2.5E-7
+ pku0 = 0 lkvth0 = 0 wkvth0 = 2E-7
+ pkvth0 = 0 stk2 = 0 lodk2 = 1
+ steta0 = 0 lodeta0 = 1

.model pshort_model.31 pmos
+ level = 54 lmin = 1.8E-7 lmax = 2.5E-7 wmin = 1E-6
+ wmax = 3E-6 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 4.23E-9
+ toxm = 4.23E-9 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 9.999999999999999E22 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {7.3039E-9+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {-1.3994E-8-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = -5.722E-9 dwb = -1.7864E-8 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = -0.898665874443435 lvth0 = -2.47045293961666E-8
+ wvth0 = -4.417326424694477E-10 pvth0 = 4.885547948940715E-15 k1 = 0.48367106012707
+ lk1 = 1.059021870017724E-7 wk1 = -1.510490758408703E-6 pk1 = 3.419975290533616E-13
+ k2 = 0.015695910369266 lk2 = -3.886777502260058E-8 wk2 = 5.586343067432635E-7
+ pk2 = -1.272034032742396E-13 k3 = -15.845 k3b = 2
+ w0 = 0 lpe0 = 0 lpeb = 0
+ vbm = -3 dvtp0 = 0 dvtp1 = 0
+ dvt0 = 4.4955 dvt1 = 0.294 dvt2 = 0.015
+ dvt0w = -4.9772 dvt1w = 1.1472E6 dvt2w = -8.96E-3
+ vfbsdoff = 0 u0 = 4.516182440855904E-3 lu0 = -1.403367379403021E-10
+ wu0 = 6.289958725098423E-9 pu0 = -1.489488917862708E-15 ua = -2.043015578595517E-9
+ lua = -2.709842405873682E-17 wua = 2.719234354385535E-15 pua = -6.070842165562616E-22
+ ub = 1.797873252787153E-18 lub = 3.84052384225212E-26 wub = -2.121175514939846E-24
+ pub = 4.819514750193827E-31 uc = -3.902944066476121E-11 luc = 8.172517531185773E-18
+ wuc = 3.800533978453389E-17 puc = -7.911753339027454E-24 ud = 0
+ up = 0 lp = 1 eu = 1.67
+ vsat = 1.704280267758007E5 lvsat = -0.015774460116019 wvsat = 0.224139640520951
+ pvsat = -4.510416641716087E-8 a0 = -0.979586871198539 la0 = 3.689372908380954E-7
+ wa0 = 9.606864420302784E-7 pa0 = -1.398127118006856E-13 ags = 0.822976281723223
+ lags = 8.88158091169503E-8 wags = -2.820150409772537E-6 pags = 5.865574434277705E-13
+ b0 = 0 b1 = 3.084995029587185E-24 lb1 = -8.575915982848829E-31
+ wb1 = -9.209920098368354E-30 pb1 = 2.560247268305222E-36 keta = -0.503714376127331
+ lketa = 1.094056916266951E-7 wketa = 3.779308792722639E-7 pketa = -7.761764947990384E-14
+ a1 = 0 a2 = 1.743083079353516 la2 = -2.243259212043906E-7
+ wa2 = -1.678973214834472E-6 pa2 = 3.537675895442328E-13 rdsw = 547.88
+ rdswmin = 0 rdw = 0 rdwmin = 0
+ rsw = 0 rswmin = 0 prwb = -0.32348
+ prwg = 0.1376 wr = 1 voff = -0.18685842374617
+ lvoff = -3.149791402635296E-8 wvoff = 1.393179668989751E-7 pvoff = -3.468168032498798E-14
+ voffl = 0 minv = 0 nfactor = 1.286512992138004
+ lnfactor = 1.420500879593939E-7 wnfactor = -7.256414746185846E-7 pnfactor = 2.222645493190001E-13
+ eta0 = 0.279640046423887 leta0 = -2.331375035938774E-8 weta0 = 1.02307646133359E-6
+ peta0 = -2.03806477050942E-13 etab = 0.301146219551655 letab = -8.372722268879616E-8
+ wetab = -2.046039838916166E-7 petab = 5.687234120048298E-14 dsub = 0.935752122700463
+ ldsub = -1.378863363910617E-7 wdsub = 7.464172682376615E-7 pdsub = -1.559245231445469E-13
+ cit = 1E-5 cdsc = 1.3E-4 cdscb = 7.8E-4
+ cdscd = 0 pclm = 1.899059771567209 lpclm = -2.628592557659633E-7
+ wpclm = -1.19927894241106E-6 ppclm = 2.467340943766432E-13 pdiblc1 = 0.812324477057923
+ lpdiblc1 = -1.284227244941422E-7 wpdiblc1 = 5.615233055025632E-7 ppdiblc1 = -1.255270065806185E-13
+ pdiblc2 = 9.927601011035878E-3 lpdiblc2 = -1.051885191858297E-9 wpdiblc2 = 2.674937616581596E-8
+ ppdiblc2 = -6.087254851238051E-15 pdiblcb = -0.408231747003947 lpdiblcb = 9.253286364543624E-8
+ wpdiblcb = -2.586229076247941E-7 ppdiblcb = 3.090506343595089E-14 drout = -0.342675617131599
+ ldrout = 2.79260416255967E-7 wdrout = -9.009153844901299E-7 pdrout = 1.873795889893332E-13
+ pscbe1 = 7.9992886E8 pscbe2 = 8.385605779847905E-9 lpscbe2 = 2.360686095721679E-16
+ wpscbe2 = 2.889198479330202E-16 ppscbe2 = -8.72022866355544E-23 pvag = 0
+ delta = 0.01 fprout = 0 pdits = 0
+ pditsl = 0 pditsd = 0 lambda = 0
+ vtl = 0 lc = 5E-9 xn = 3
+ alpha0 = 1E-10 alpha1 = 1E-10 beta0 = 9.52359642714142
+ lbeta0 = -2.178170346211925E-7 wbeta0 = 1.239177095039083E-6 pbeta0 = -1.929631678173612E-13
+ aigbacc = 0.43 bigbacc = 0.054 cigbacc = 0.075
+ nigbacc = 1 aigbinv = 0.35 bigbinv = 0.03
+ cigbinv = 6E-3 eigbinv = 1.1 nigbinv = 3
+ aigc = 0.43 bigc = 0.054 cigc = 0.075
+ aigsd = 0.43 bigsd = 0.054 cigsd = 0.075
+ dlcig = 0 nigc = 1 poxedge = 1
+ pigcd = 1 ntox = 1 toxref = 4.23E-9
+ agidl = 1.380571860329356E-8 lagidl = -2.788044899508319E-15 wagidl = -1.350550820708037E-14
+ pagidl = 2.747317697225282E-21 bgidl = 4.616408933089225E8 lbgidl = 111.66958458236586
+ wbgidl = 1.607213077914511E3 pbgidl = -3.333775067894354E-4 cgidl = -1.118076363127147E3
+ lcgidl = 2.94942866614089E-4 wcgidl = 1.397361387229858E-3 pcgidl = -2.906344002071637E-10
+ egidl = 7.603999023644048 legidl = -1.560741748929679E-6 wegidl = -7.394382106706462E-6
+ pegidl = 1.537942745609664E-12 noia = 1.5E42 noib = 0
+ noic = 0 em = 4.1E7 af = 1
+ ef = 1 kf = 0 lintnoi = -2E-7
+ tnoia = 2.5E7 tnoib = 0 ntnoi = 1
+ rnoia = 0.69 rnoib = 0.34 xpart = 0
+ cgso = {5.248925E-11/sw_func_tox_lv_ratio} cgdo = {5.248925E-11/sw_func_tox_lv_ratio} cgbo = {0/sw_func_tox_lv_ratio}
+ ckappas = 0.6 cf = 1.2E-11 clc = 1E-7
+ cle = 0.6 dlc = -3E-9 dwc = 0
+ vfbcv = -0.14469 noff = 3.9 voffcv = -0.10701
+ acde = 0.8 moin = 18.13 cgsl = {9.548271750000001E-12/sw_func_tox_lv_ratio}
+ cgdl = {9.548271750000001E-12/sw_func_tox_lv_ratio} ijthsrev = 0.1 ijthsfwd = 0.1
+ xjbvs = 1 bvs = 12.69 jss = 2.1483E-5
+ jsws = 8.040000000000001E-10 cjs = {sw_psd_nw_cj} mjs = 0.34629
+ mjsws = 0.29781 cjsws = {9.888891999999999E-11*sw_func_psd_nw_cj} cjswgs = {2.39155046E-10*sw_func_psd_nw_cj}
+ mjswgs = 0.9274 pbs = 0.6587 pbsws = 0.7418
+ pbswgs = 1.4338 xrcrg1 = 12 xrcrg2 = 1
+ rbpb = 50 rbpd = 50 rbps = 50
+ rbdb = 50 rbsb = 50 gbmin = 1E-12
+ tnom = 30 ute = -0.401747722602166 lute = 1.257081168727968E-8
+ wute = 3.037568574242714E-7 pute = -3.752880315887361E-14 kt1 = -0.4465487668033
+ lkt1 = -2.739284604212753E-8 wkt1 = 3.04374721618198E-7 pkt1 = -7.556787168928261E-14
+ kt1l = 0 kt2 = 0.038929515336004 lkt2 = -3.36639392735405E-8
+ wkt2 = 2.441397724318327E-7 pkt2 = -5.017852470274515E-14 ua1 = 3.2654354721609E-11
+ lua1 = 1.95803295921868E-17 wua1 = 1.102418654310764E-15 pua1 = -2.244317192469641E-22
+ ub1 = 3.6988817057E-19 wub1 = 6.810225764805252E-26 uc1 = 1.154503318194338E-12
+ luc1 = -1.501701269253182E-19 wuc1 = -1.654066454521496E-18 puc1 = 4.483167255958548E-25
+ at = -1.344075929300765E4 lat = 0.017944634881481 wat = 0.100529433610427
+ pat = -2.371519060088096E-8 prt = 0 njs = 1.3632
+ xtis = 5.2 tpb = 2.0386E-3 tpbsw = 1.246E-3
+ tpbswg = 0 tcj = 1.2407E-3 tcjsw = 3.7357E-4
+ tcjswg = 2E-12 tvoff = 0 tvfbsdoff = 0
+ saref = 1.25E-6 sbref = 1.24E-6 wlod = 0
+ ku0 = 4.5E-8 kvsat = 0.5 kvth0 = 3.29E-8
+ tku0 = 0 llodku0 = 0 wlodku0 = 1
+ llodvth = 0 wlodvth = 1 lku0 = 0
+ wku0 = 2.5E-7 pku0 = 0 lkvth0 = 0
+ wkvth0 = 2E-7 pkvth0 = 0 stk2 = 0
+ lodk2 = 1 steta0 = 0 lodeta0 = 1

.model pshort_model.32 pmos
+ level = 54 lmin = 1.5E-7 lmax = 1.8E-7 wmin = 1E-6
+ wmax = 3E-6 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 4.23E-9
+ toxm = 4.23E-9 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 9.999999999999999E22 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {7.3039E-9+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {-1.3994E-8-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = -5.722E-9 dwb = -1.7864E-8 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = -0.804969765443255 lvth0 = -4.419219571489606E-8
+ wvth0 = 2.210796835696688E-8 pvth0 = 1.954807374699516E-16 k1 = -0.401689142682068
+ lk1 = 2.900464848636393E-7 wk1 = -6.480368568297199E-7 pk1 = 1.62617466971752E-13
+ k2 = 0.428132653805264 lk2 = -1.24649668416367E-7 wk2 = 1.944470702032923E-7
+ pk2 = -5.145682832076403E-14 k3 = -15.845 k3b = 2
+ w0 = 0 lpe0 = 0 lpeb = 0
+ vbm = -3 dvtp0 = 0 dvtp1 = 0
+ dvt0 = 4.4955 dvt1 = 0.294 dvt2 = 0.015
+ dvt0w = -4.9772 dvt1w = 1.1472E6 dvt2w = -8.96E-3
+ vfbsdoff = 0 u0 = 6.784521537583039E-3 lu0 = -6.121240499903856E-10
+ wu0 = -1.328912397545169E-9 pu0 = 9.514484919368745E-17 ua = -6.699130238097632E-10
+ lua = -3.126872782235161E-16 wua = -4.065997816336757E-16 pua = 4.305177372610201E-23
+ ub = 4.754108914380993E-19 lub = 3.134615400347882E-25 wub = 3.711512341085188E-25
+ pub = -3.64225808616886E-32 uc = 7.623933468844942E-13 luc = -1.037064412283932E-19
+ wuc = -5.425409594631171E-19 puc = 1.057432811549956E-25 ud = 0
+ up = 0 lp = 1 eu = 1.67
+ vsat = 3.262428220498732E5 lvsat = -0.048182067755482 wvsat = 0.051018477125728
+ pvsat = -9.097041884915179E-9 a0 = 0.102571675072607 la0 = 1.438612991162522E-7
+ wa0 = 3.080820608533956E-6 pa0 = -5.807751768234525E-13 ags = 1.25
+ b0 = 0 b1 = -7.198321735703424E-24 lb1 = 1.281214889094382E-30
+ wb1 = 2.148981356285948E-29 pb1 = -3.824928936426233E-36 keta = 0.027382427553184
+ lketa = -1.056070377207871E-9 wketa = 1.605140337412628E-7 pketa = -3.239755461160198E-14
+ a1 = 0 a2 = -1.322818789860381 la2 = 4.133448767696694E-7
+ wa2 = 1.520436179080246E-7 pa2 = -2.706193946421349E-14 rdsw = 547.88
+ rdswmin = 0 rdw = 0 rdwmin = 0
+ rsw = 0 rswmin = 0 prwb = -0.32348
+ prwg = 0.1376 wr = 1 voff = 0.010515769173285
+ lvoff = -7.254937766328454E-8 wvoff = -2.558120482846986E-7 pvoff = 4.750062127303394E-14
+ voffl = 0 minv = 0 nfactor = -2.655313189523576
+ lnfactor = 9.619026318308228E-7 wnfactor = 2.458026897902803E-6 pnfactor = -4.399002681449782E-13
+ eta0 = -0.767055570458474 leta0 = 1.943863776047408E-7 weta0 = 1.986469742676889E-7
+ peta0 = -3.233503689507946E-14 etab = -0.580051309957149 letab = 9.955128907868101E-8
+ wetab = 3.560066669517047E-7 petab = -5.972794684711775E-14 dsub = 0.367115443023737
+ ldsub = -1.961673065845884E-8 wdsub = -7.750113975429845E-8 pdsub = 1.544061869688482E-14
+ cit = 1E-5 cdsc = 1.3E-4 cdscb = 7.8E-4
+ cdscd = 0 pclm = 1.803740738075466 lpclm = -2.430340406280826E-7
+ wpclm = -1.804094770424366E-7 ppclm = 3.482147201355395E-14 pdiblc1 = 1.235341761339374
+ lpdiblc1 = -2.164052434172724E-7 wpdiblc1 = -2.912299105250456E-7 ppdiblc1 = 5.183542931453181E-14
+ pdiblc2 = 0.031213394907501 lpdiblc2 = -5.4790748927963E-9 wpdiblc2 = -1.745685337541072E-8
+ ppdiblc2 = 3.107110418582602E-15 pdiblcb = 0.254544669229239 lpdiblcb = -4.531667761407183E-8
+ wpdiblcb = -7.630579827320235E-7 ppdiblcb = 1.358215058373533E-13 drout = 1
+ pscbe1 = 8E8 pscbe2 = 8.761485201233655E-9 lpscbe2 = 1.578902004769882E-16
+ wpscbe2 = 6.890437900600571E-16 ppscbe2 = -1.704232651106726E-22 pvag = 0
+ delta = 0.01 fprout = 0 pdits = 0
+ pditsl = 0 pditsd = 0 lambda = 0
+ vtl = 0 lc = 5E-9 xn = 3
+ alpha0 = 1E-10 alpha1 = 1E-10 beta0 = 14.58396122072988
+ lbeta0 = -1.270312187310069E-6 wbeta0 = 3.302930127020686E-6 pbeta0 = -6.22199033433151E-13
+ aigbacc = 0.43 bigbacc = 0.054 cigbacc = 0.075
+ nigbacc = 1 aigbinv = 0.35 bigbinv = 0.03
+ cigbinv = 6E-3 eigbinv = 1.1 nigbinv = 3
+ aigc = 0.43 bigc = 0.054 cigc = 0.075
+ aigsd = 0.43 bigsd = 0.054 cigsd = 0.075
+ dlcig = 0 nigc = 1 poxedge = 1
+ pigcd = 1 ntox = 1 toxref = 4.23E-9
+ agidl = 3.063054396323376E-9 lagidl = -5.536996564290045E-16 wagidl = -7.713078303536958E-15
+ pagidl = 1.542561786447095E-21 bgidl = 9.899116899967341E8 lbgidl = 1.795598120861303
+ wbgidl = 30.11756199493219 pbgidl = -5.36056462435399E-6 cgidl = 300
+ egidl = 0.1 noia = 1.5E42 noib = 0
+ noic = 0 em = 4.1E7 af = 1
+ ef = 1 kf = 0 lintnoi = -2E-7
+ tnoia = 2.5E7 tnoib = 0 ntnoi = 1
+ rnoia = 0.69 rnoib = 0.34 xpart = 0
+ cgso = {5.248925E-11/sw_func_tox_lv_ratio} cgdo = {5.248925E-11/sw_func_tox_lv_ratio} cgbo = {0/sw_func_tox_lv_ratio}
+ ckappas = 0.6 cf = 1.2E-11 clc = 1E-7
+ cle = 0.6 dlc = -3E-9 dwc = 0
+ vfbcv = -0.14469 noff = 3.9 voffcv = -0.10701
+ acde = 0.8 moin = 18.13 cgsl = {9.548271750000001E-12/sw_func_tox_lv_ratio}
+ cgdl = {9.548271750000001E-12/sw_func_tox_lv_ratio} ijthsrev = 0.1 ijthsfwd = 0.1
+ xjbvs = 1 bvs = 12.69 jss = 2.1483E-5
+ jsws = 8.040000000000001E-10 cjs = {sw_psd_nw_cj} mjs = 0.34629
+ mjsws = 0.29781 cjsws = {9.888891999999999E-11*sw_func_psd_nw_cj} cjswgs = {2.39155046E-10*sw_func_psd_nw_cj}
+ mjswgs = 0.9274 pbs = 0.6587 pbsws = 0.7418
+ pbswgs = 1.4338 xrcrg1 = 12 xrcrg2 = 1
+ rbpb = 50 rbpd = 50 rbps = 50
+ rbdb = 50 rbsb = 50 gbmin = 1E-12
+ tnom = 30 ute = -0.330404354505448 lute = -2.267752756420609E-9
+ wute = 9.07689227865991E-8 pute = 6.770131390546588E-15 kt1 = 0.071255523490432
+ lkt1 = -1.350899247717402E-7 wkt1 = -2.799133286792807E-7 pkt1 = 4.595703131598939E-14
+ kt1l = 0 kt2 = -0.122925684356 wkt2 = 2.882946544064429E-9
+ ua1 = 1.452037965373941E-12 lua1 = 2.607003704968262E-17 wua1 = 3.975585951480688E-16
+ pua1 = -7.78292852618335E-23 ub1 = 1.650057705471264E-19 lub1 = 4.261308061595746E-26
+ wub1 = 6.797565765936195E-25 pub1 = -1.272167584888506E-31 uc1 = -3.101281976675811E-10
+ luc1 = 6.459289628570414E-17 wuc1 = 2.654867631892407E-16 puc1 = -5.511377015035095E-23
+ at = 2.301444998112198E5 lat = -0.032718175989089 wat = 0.053860177339858
+ pat = -1.400854532767796E-8 prt = 0 njs = 1.3632
+ xtis = 5.2 tpb = 2.0386E-3 tpbsw = 1.246E-3
+ tpbswg = 0 tcj = 1.2407E-3 tcjsw = 3.7357E-4
+ tcjswg = 2E-12 tvoff = 0 tvfbsdoff = 0
+ saref = 1.1E-6 sbref = 1.1E-6 wlod = 0
+ ku0 = 4.5E-8 kvsat = 0.5 kvth0 = 3.29E-8
+ tku0 = 0 llodku0 = 0 wlodku0 = 1
+ llodvth = 0 wlodvth = 1 lku0 = 0
+ wku0 = 2.5E-7 pku0 = 0 lkvth0 = 0
+ wkvth0 = 2E-7 pkvth0 = 0 stk2 = 0
+ lodk2 = 1 steta0 = 0 lodeta0 = 1

.model pshort_model.33 pmos
+ level = 54 lmin = 8E-6 lmax = 2.02E-5 wmin = 5.5E-7
+ wmax = 1E-6 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 4.23E-9
+ toxm = 4.23E-9 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 9.999999999999999E22 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {7.3039E-9+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {-1.3994E-8-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = -5.722E-9 dwb = -1.7864E-8 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = -0.993400837766711 wvth0 = -2.598101060861724E-8
+ k1 = 0.507360724147231 wk1 = -1.536295825918915E-8 k2 = -3.335314292170001E-3
+ wk2 = 6.356442781794394E-10 k3 = -15.845 k3b = 2
+ w0 = 0 lpe0 = 0 lpeb = 0
+ vbm = -3 dvtp0 = 0 dvtp1 = 0
+ dvt0 = 4.4955 dvt1 = 0.294 dvt2 = 0.015
+ dvt0w = -4.9772 dvt1w = 1.1472E6 dvt2w = -8.96E-3
+ vfbsdoff = 0 u0 = 3.576710462304844E-3 wu0 = 2.616329352629852E-9
+ ua = -2.003411319904672E-9 wua = 5.831326566317479E-16 ub = 1.787490124338378E-18
+ wub = -4.113008560176676E-25 uc = -4.302947739237318E-12 wuc = -3.410801900969911E-17
+ ud = 0 up = 0 lp = 1
+ eu = 1.67 vsat = 9.181913986396312E4 wvsat = -0.036046950215831
+ a0 = 1.1662826684512 wa0 = 4.53204847680015E-8 ags = 0.351217706664413
+ wags = -6.224184174572695E-8 b0 = 8.948902158933335E-8 wb0 = -8.818178385976069E-14
+ b1 = 1.540739775555556E-11 wb1 = -1.518232957062195E-17 keta = 5.727252612387334E-3
+ wketa = 8.996479898929582E-10 a1 = 0 a2 = 0.8
+ rdsw = 547.88 rdswmin = 0 rdw = 0
+ rdwmin = 0 rsw = 0 rswmin = 0
+ prwb = -0.32348 prwg = 0.1376 wr = 1
+ voff = -0.209936786628644 wvoff = -4.189801252097148E-8 voffl = 0
+ minv = 0 nfactor = 1.444085569201378 wnfactor = 1.131498575765622E-7
+ eta0 = 0.08 etab = -0.07 dsub = 0.56
+ cit = 1E-5 cdsc = 1.3E-4 cdscb = 7.8E-4
+ cdscd = 0 pclm = 1.7402344E-3 pdiblc1 = 0.39
+ pdiblc2 = 2.465593676892934E-4 wpdiblc2 = 3.165857933389863E-10 pdiblcb = -0.225
+ drout = 0.56 pscbe1 = 8.117496174794577E8 wpscbe1 = -11.592476536503357
+ pscbe2 = 1.226411215477716E-8 wpscbe2 = -1.470344255216402E-15 pvag = 0
+ delta = 0.01 fprout = 0 pdits = 0
+ pditsl = 0 pditsd = 0 lambda = 0
+ vtl = 0 lc = 5E-9 xn = 3
+ alpha0 = -1.189760444444445E-10 walpha0 = 1.172380661824089E-16 alpha1 = -1.189760444444445E-10
+ walpha1 = 1.172380661824089E-16 beta0 = 62.12353200000001 wbeta0 = -3.165427786925041E-5
+ aigbacc = 0.43 bigbacc = 0.054 cigbacc = 0.075
+ nigbacc = 1 aigbinv = 0.35 bigbinv = 0.03
+ cigbinv = 6E-3 eigbinv = 1.1 nigbinv = 3
+ aigc = 0.43 bigc = 0.054 cigc = 0.075
+ aigsd = 0.43 bigsd = 0.054 cigsd = 0.075
+ dlcig = 0 nigc = 1 poxedge = 1
+ pigcd = 1 ntox = 1 toxref = 4.23E-9
+ agidl = -1.074532685381716E-9 wagidl = 1.203400986574265E-15 bgidl = 1E9
+ cgidl = 300 egidl = 0.1 noia = 1.5E42
+ noib = 0 noic = 0 em = 4.1E7
+ af = 1 ef = 1 kf = 0
+ lintnoi = -2E-7 tnoia = 2.5E7 tnoib = 0
+ ntnoi = 1 rnoia = 0.69 rnoib = 0.34
+ xpart = 0 cgso = {5.248925E-11/sw_func_tox_lv_ratio} cgdo = {5.248925E-11/sw_func_tox_lv_ratio}
+ cgbo = {0/sw_func_tox_lv_ratio} ckappas = 0.6 cf = 1.2E-11
+ clc = 1E-7 cle = 0.6 dlc = -3E-9
+ dwc = 0 vfbcv = -0.14469 noff = 3.9
+ voffcv = -0.10701 acde = 0.8 moin = 18.13
+ cgsl = {9.548271750000001E-12/sw_func_tox_lv_ratio} cgdl = {9.548271750000001E-12/sw_func_tox_lv_ratio} ijthsrev = 0.1
+ ijthsfwd = 0.1 xjbvs = 1 bvs = 12.69
+ jss = 2.1483E-5 jsws = 8.040000000000001E-10 cjs = {sw_psd_nw_cj}
+ mjs = 0.34629 mjsws = 0.29781 cjsws = {9.888891999999999E-11*sw_func_psd_nw_cj}
+ cjswgs = {2.39155046E-10*sw_func_psd_nw_cj} mjswgs = 0.9274 pbs = 0.6587
+ pbsws = 0.7418 pbswgs = 1.4338 xrcrg1 = 12
+ xrcrg2 = 1 rbpb = 50 rbpd = 50
+ rbps = 50 rbdb = 50 rbsb = 50
+ gbmin = 1E-12 tnom = 30 ute = -1.2595
+ kt1 = -0.569405208888889 wkt1 = 2.34476132364818E-8 kt1l = 0
+ kt2 = -0.052484 ua1 = -2.5605E-10 ub1 = 4.9434E-19
+ uc1 = 8.1951E-12 at = 1E4 prt = 0
+ njs = 1.3632 xtis = 5.2 tpb = 2.0386E-3
+ tpbsw = 1.246E-3 tpbswg = 0 tcj = 1.2407E-3
+ tcjsw = 3.7357E-4 tcjswg = 2E-12 tvoff = 0
+ tvfbsdoff = 0 saref = 3E-6 sbref = 3E-6
+ wlod = 0 ku0 = 4.5E-8 kvsat = 0.5
+ kvth0 = 3.29E-8 tku0 = 0 llodku0 = 0
+ wlodku0 = 1 llodvth = 0 wlodvth = 1
+ lku0 = 0 wku0 = 2.5E-7 pku0 = 0
+ lkvth0 = 0 wkvth0 = 2E-7 pkvth0 = 0
+ stk2 = 0 lodk2 = 1 steta0 = 0
+ lodeta0 = 1

.model pshort_model.34 pmos
+ level = 54 lmin = 4E-6 lmax = 8E-6 wmin = 5.5E-7
+ wmax = 1E-6 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 4.23E-9
+ toxm = 4.23E-9 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 9.999999999999999E22 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {7.3039E-9+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {-1.3994E-8-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = -5.722E-9 dwb = -1.7864E-8 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = -0.944039522207394 lvth0 = -3.962720489744132E-7
+ wvth0 = -7.137847206172534E-8 pvth0 = 3.644502757760143E-13 k1 = 0.58049642306484
+ lk1 = -5.871325132821761E-7 wk1 = -4.574285058926025E-8 pk1 = 2.438894110671028E-13
+ k2 = -9.852573571886831E-3 lk2 = 5.232047929045536E-8 wk2 = -4.934909140601843E-9
+ pk2 = 4.47203359993351E-14 k3 = -15.845 k3b = 2
+ w0 = 0 lpe0 = 0 lpeb = 0
+ vbm = -3 dvtp0 = 0 dvtp1 = 0
+ dvt0 = 4.4955 dvt1 = 0.294 dvt2 = 0.015
+ dvt0w = -4.9772 dvt1w = 1.1472E6 dvt2w = -8.96E-3
+ vfbsdoff = 0 u0 = -3.082385649855187E-3 lu0 = 5.345914367926738E-8
+ wu0 = 6.983336134771561E-9 pu0 = -3.505827804295225E-14 ua = -3.195320923830041E-9
+ lua = 9.568635997397616E-15 wua = 1.185250020685244E-15 pua = -4.833790973213096E-21
+ ub = 2.137688986406309E-18 lub = -2.811392262295012E-24 wub = -3.735036389537853E-25
+ pub = -3.034356050222422E-31 uc = 2.46171558385188E-11 luc = -2.321702444809832E-16
+ wuc = -4.707237816193425E-17 puc = 1.040777197018338E-22 ud = 0
+ up = 0 lp = 1 eu = 1.67
+ vsat = 1.570856207444297E5 lvsat = -0.523958525310615 wvsat = -0.087964335690025
+ pvsat = 4.167921475782012E-7 a0 = 1.333039775391511 la0 = -1.338724053431532E-6
+ wa0 = -4.235840523190971E-8 pa0 = 7.038850767726072E-13 ags = 0.231741355247949
+ lags = 9.591547154551625E-7 wags = 2.221977392788216E-9 pags = -5.1751476647817E-13
+ b0 = 1.99866214735941E-7 lb0 = -8.861067820546481E-13 wb0 = -1.969466090443213E-13
+ pb0 = 8.731627114037501E-19 b1 = 2.14636985376576E-10 lb1 = -1.599412738666501E-15
+ wb1 = -2.115016112215921E-16 pb1 = 1.576048837262608E-21 keta = 0.017135704001098
+ lketa = -9.15869108471508E-8 wketa = -6.950667897939236E-9 pketa = 6.302224174372618E-14
+ a1 = 0 a2 = 0.8 rdsw = 547.88
+ rdswmin = 0 rdw = 0 rdwmin = 0
+ rsw = 0 rswmin = 0 prwb = -0.32348
+ prwg = 0.1376 wr = 1 voff = -0.162560385566834
+ lvoff = -3.803371792073992E-7 wvoff = -9.974985397703775E-8 pvoff = 4.644338889872025E-13
+ voffl = 0 minv = 0 nfactor = 0.876308540435568
+ lnfactor = 4.558107173607574E-6 wnfactor = 2.694436882819492E-7 pnfactor = -1.254724997376879E-12
+ eta0 = 0.08 etab = -0.07 dsub = 0.56
+ cit = 1E-5 cdsc = 1.3E-4 cdscb = 7.8E-4
+ cdscd = 0 pclm = 0.398721529855687 lpclm = -3.186961076142708E-6
+ wpclm = -4.271659716960183E-7 ppclm = 3.429283294783974E-12 pdiblc1 = 0.39
+ pdiblc2 = -1.278604057430475E-3 lpdiblc2 = 1.22439936749004E-8 wpdiblc2 = 1.353047461158289E-9
+ ppdiblc2 = -8.320701831713345E-15 pdiblcb = -0.225 drout = 0.56
+ pscbe1 = 8.235814911340632E8 lpscbe1 = -94.98613971668921 wpscbe1 = -23.266089243008818
+ ppscbe1 = 9.371562272447334E-5 pscbe2 = 1.513626549107818E-8 lpscbe2 = -2.305761251798459E-14
+ wpscbe2 = -3.041239461028293E-15 ppscbe2 = 1.261112786151539E-20 pvag = 0
+ delta = 0.01 fprout = 0 pdits = 0
+ pditsl = 0 pditsd = 0 lambda = 0
+ vtl = 0 lc = 5E-9 xn = 3
+ alpha0 = -2.132866011838728E-10 lalpha0 = 7.571240177774496E-16 walpha0 = 2.10170953171099E-16
+ palpha0 = -7.460641015505601E-22 alpha1 = -2.387845239880348E-10 lalpha1 = 9.618210360741879E-16
+ walpha1 = 2.352964074185223E-16 palpha1 = -9.477709467434233E-22 beta0 = 86.88298219284056
+ lbeta0 = -1.987685690347216E-4 wbeta0 = -5.605204696556397E-5 pbeta0 = 1.958649975319762E-10
+ aigbacc = 0.43 bigbacc = 0.054 cigbacc = 0.075
+ nigbacc = 1 aigbinv = 0.35 bigbinv = 0.03
+ cigbinv = 6E-3 eigbinv = 1.1 nigbinv = 3
+ aigc = 0.43 bigc = 0.054 cigc = 0.075
+ aigsd = 0.43 bigsd = 0.054 cigsd = 0.075
+ dlcig = 0 nigc = 1 poxedge = 1
+ pigcd = 1 ntox = 1 toxref = 4.23E-9
+ agidl = -2.38402859155395E-9 lagidl = 1.051261742079983E-14 wagidl = 2.483080462587838E-15
+ pagidl = -1.027325147728325E-20 bgidl = 1.385342418682815E9 lbgidl = -3.093524313076614E3
+ wbgidl = -379.71341369918014 pbgidl = 3.048334728616054E-3 cgidl = 300
+ egidl = 0.1 noia = 1.5E42 noib = 0
+ noic = 0 em = 4.1E7 af = 1
+ ef = 1 kf = 0 lintnoi = -2E-7
+ tnoia = 2.5E7 tnoib = 0 ntnoi = 1
+ rnoia = 0.69 rnoib = 0.34 xpart = 0
+ cgso = {5.248925E-11/sw_func_tox_lv_ratio} cgdo = {5.248925E-11/sw_func_tox_lv_ratio} cgbo = {0/sw_func_tox_lv_ratio}
+ ckappas = 0.6 cf = 1.2E-11 clc = 1E-7
+ cle = 0.6 dlc = -3E-9 dwc = 0
+ vfbcv = -0.14469 noff = 3.9 voffcv = -0.10701
+ acde = 0.8 moin = 18.13 cgsl = {9.548271750000001E-12/sw_func_tox_lv_ratio}
+ cgdl = {9.548271750000001E-12/sw_func_tox_lv_ratio} ijthsrev = 0.1 ijthsfwd = 0.1
+ xjbvs = 1 bvs = 12.69 jss = 2.1483E-5
+ jsws = 8.040000000000001E-10 cjs = {sw_psd_nw_cj} mjs = 0.34629
+ mjsws = 0.29781 cjsws = {9.888891999999999E-11*sw_func_psd_nw_cj} cjswgs = {2.39155046E-10*sw_func_psd_nw_cj}
+ mjswgs = 0.9274 pbs = 0.6587 pbsws = 0.7418
+ pbswgs = 1.4338 xrcrg1 = 12 xrcrg2 = 1
+ rbpb = 50 rbpd = 50 rbps = 50
+ rbdb = 50 rbsb = 50 gbmin = 1E-12
+ tnom = 30 ute = -2.809380267012881 lute = 1.24424201850162E-5
+ wute = 3.469145523671752E-7 pute = -2.785025863429054E-12 kt1 = -0.596421808266296
+ lkt1 = 2.168889356026298E-7 wkt1 = -3.361000226770598E-8 pkt1 = 4.580578525762334E-13
+ kt1l = 0 kt2 = -0.116488052725888 lkt2 = 5.13823767234798E-7
+ wkt2 = 3.752564264789023E-8 pkt2 = -3.01255408869551E-13 ua1 = -4.297832865011864E-9
+ lua1 = 3.244738433892087E-14 wua1 = 1.823872121172453E-15 pua1 = -1.4642023502307E-20
+ ub1 = 3.738579573427357E-18 lub1 = -2.604471636459993E-23 wub1 = -1.698653782777586E-24
+ pub1 = 1.363677218429306E-29 uc1 = 1.396602447982411E-10 luc1 = -1.055400604858542E-15
+ wuc1 = -4.20298780128007E-17 puc1 = 3.374153563282278E-22 at = -2.656065136339185E4
+ lat = 0.293508470417493 wat = -8.892762891253798E-3 pat = 7.139099377783079E-8
+ prt = 0 njs = 1.3632 xtis = 5.2
+ tpb = 2.0386E-3 tpbsw = 1.246E-3 tpbswg = 0
+ tcj = 1.2407E-3 tcjsw = 3.7357E-4 tcjswg = 2E-12
+ tvoff = 0 tvfbsdoff = 0 saref = 3E-6
+ sbref = 3E-6 wlod = 0 ku0 = 4.5E-8
+ kvsat = 0.5 kvth0 = 3.29E-8 tku0 = 0
+ llodku0 = 0 wlodku0 = 1 llodvth = 0
+ wlodvth = 1 lku0 = 0 wku0 = 2.5E-7
+ pku0 = 0 lkvth0 = 0 wkvth0 = 2E-7
+ pkvth0 = 0 stk2 = 0 lodk2 = 1
+ steta0 = 0 lodeta0 = 1

.model pshort_model.35 pmos
+ level = 54 lmin = 2E-6 lmax = 4E-6 wmin = 5.5E-7
+ wmax = 1E-6 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 4.23E-9
+ toxm = 4.23E-9 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 9.999999999999999E22 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {7.3039E-9+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {-1.3994E-8-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = -5.722E-9 dwb = -1.7864E-8 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = -1.094543031462421 lvth0 = 2.099542802627264E-7
+ wvth0 = 6.745391093192534E-8 pvth0 = -1.947648969338147E-13 k1 = 0.393618983351444
+ lk1 = 1.656075713541076E-7 wk1 = 4.385127259054034E-8 pk1 = -1.169946419716561E-13
+ k2 = 3.632959699180497E-3 lk2 = -1.999086899004571E-9 wk2 = 9.167005326286113E-9
+ pk2 = -1.208200625031599E-14 k3 = -15.845 k3b = 2
+ w0 = 0 lpe0 = 0 lpeb = 0
+ vbm = -3 dvtp0 = 0 dvtp1 = 0
+ dvt0 = 4.4955 dvt1 = 0.294 dvt2 = 0.015
+ dvt0w = -4.9772 dvt1w = 1.1472E6 dvt2w = -8.96E-3
+ vfbsdoff = 0 u0 = 0.015234805161733 lu0 = -2.032228110352153E-8
+ wu0 = -6.085898307123801E-9 pu0 = 1.758444145818896E-14 ua = -1.278216710812904E-10
+ lua = -2.787214182683316E-15 wua = -5.023687525516261E-16 pua = 1.963917193959736E-21
+ ub = 1.46065485336248E-18 lub = -8.430689880406223E-26 wub = -6.277719535075555E-25
+ pub = 7.207541147805693E-31 uc = -4.664542664722006E-11 luc = 5.487458262058315E-17
+ wuc = -1.73398932781645E-17 puc = -1.568437262017212E-23 ud = 0
+ up = 0 lp = 1 eu = 1.67
+ vsat = -2.530485752884978E4 lvsat = 0.210708132488415 wvsat = 0.056373575775961
+ pvsat = -1.645992277518505E-7 a0 = 1.063759530135458 la0 = -2.540664569030965E-7
+ wa0 = 1.45395715396801E-7 pa0 = -5.238626807039213E-14 ags = 0.654870180860539
+ lags = -7.452031165664424E-7 wags = -4.080978973563052E-7 pags = 1.135248765172681E-12
+ b0 = -1.306126969197936E-7 lb0 = 4.450583083477107E-13 wb0 = 1.287047327657286E-13
+ pb0 = -4.38556985591029E-19 b1 = -9.122121007252772E-11 lb1 = -3.674195976958562E-16
+ wb1 = 8.988866888003025E-17 pb1 = 3.620524056966348E-22 keta = -6.992750127050394E-3
+ lketa = 5.602212839580494E-9 wketa = 1.80959625365876E-8 pketa = -3.786528508698268E-14
+ a1 = 0 a2 = 0.8 rdsw = 547.88
+ rdswmin = 0 rdw = 0 rdwmin = 0
+ rsw = 0 rswmin = 0 prwb = -0.32348
+ prwg = 0.1376 wr = 1 voff = -0.288882124831054
+ lvoff = 1.284852706880061E-7 wvoff = 5.024613593888214E-8 pvoff = -1.397481584422439E-13
+ voffl = 0 minv = 0 nfactor = 2.766201122471184
+ lnfactor = -3.054357468120902E-6 wnfactor = -4.867762894389234E-7 pnfactor = 1.791319998243063E-12
+ eta0 = 0.160612523 leta0 = -3.24706275293724E-7 etab = -0.140472579691598
+ letab = 2.838627053268009E-7 petab = 7.134745191146275E-21 dsub = 0.8641982
+ ldsub = -1.2253066992216E-6 cit = 1E-5 cdsc = 1.3E-4
+ cdscb = 7.8E-4 cdscd = 0 pclm = -1.209948579794565
+ lpclm = 3.292742821487189E-6 wpclm = 9.15695735221605E-7 ppclm = -1.979747546339729E-12
+ pdiblc1 = 0.39 pdiblc2 = 3.418039535498608E-3 lpdiblc2 = -6.674030357694831E-9
+ wpdiblc2 = -1.523171436371584E-9 ppdiblc2 = 3.264673372910211E-15 pdiblcb = 0.0162819904208
+ lpdiblcb = -9.718809620310977E-7 wpdiblcb = -2.377573913611311E-7 ppdiblcb = 9.576839193139397E-13
+ drout = 0.56 pscbe1 = 8E8 pscbe2 = 9.640534824161437E-9
+ lpscbe2 = -9.208753404119522E-16 wpscbe2 = -5.004272546917018E-18 ppscbe2 = 3.8120895713467E-22
+ pvag = 0 delta = 0.01 fprout = 0
+ pdits = 0 pditsl = 0 pditsd = 0
+ lambda = 0 vtl = 0 lc = 5E-9
+ xn = 3 alpha0 = -5.328414943259614E-11 lalpha0 = 1.126360621527282E-16
+ walpha0 = 4.945929298139349E-17 palpha0 = -9.871946284634858E-23 alpha1 = 5.798452524893272E-15
+ lalpha1 = -2.351723251700458E-20 walpha1 = -2.792281755779786E-21 palpha1 = 1.140605890041792E-26
+ beta0 = 72.55553832112695 lbeta0 = -1.410577970487856E-4 wbeta0 = -1.495598751037598E-5
+ pbeta0 = 3.033056319919236E-11 aigbacc = 0.43 bigbacc = 0.054
+ cigbacc = 0.075 nigbacc = 1 aigbinv = 0.35
+ bigbinv = 0.03 cigbinv = 6E-3 eigbinv = 1.1
+ nigbinv = 3 aigc = 0.43 bigc = 0.054
+ cigc = 0.075 aigsd = 0.43 bigsd = 0.054
+ cigsd = 0.075 dlcig = 0 nigc = 1
+ poxedge = 1 pigcd = 1 ntox = 1
+ toxref = 4.23E-9 agidl = 3.279837269670886E-10 lagidl = -4.113356540550982E-16
+ wagidl = -2.588439225215974E-16 pagidl = 7.711870428449332E-22 bgidl = 2.293151626343703E8
+ lbgidl = 1.562939601959449E3 wbgidl = 759.42682739836 pbgidl = -1.540108492841946E-3
+ cgidl = 300 egidl = 0.1 noia = 1.5E42
+ noib = 0 noic = 0 em = 4.1E7
+ af = 1 ef = 1 kf = 0
+ lintnoi = -2E-7 tnoia = 2.5E7 tnoib = 0
+ ntnoi = 1 rnoia = 0.69 rnoib = 0.34
+ xpart = 0 cgso = {5.248925E-11/sw_func_tox_lv_ratio} cgdo = {5.248925E-11/sw_func_tox_lv_ratio}
+ cgbo = {0/sw_func_tox_lv_ratio} ckappas = 0.6 cf = 1.2E-11
+ clc = 1E-7 cle = 0.6 dlc = -3E-9
+ dwc = 0 vfbcv = -0.14469 noff = 3.9
+ voffcv = -0.10701 acde = 0.8 moin = 18.13
+ cgsl = {9.548271750000001E-12/sw_func_tox_lv_ratio} cgdl = {9.548271750000001E-12/sw_func_tox_lv_ratio} ijthsrev = 0.1
+ ijthsfwd = 0.1 xjbvs = 1 bvs = 12.69
+ jss = 2.1483E-5 jsws = 8.040000000000001E-10 cjs = {sw_psd_nw_cj}
+ mjs = 0.34629 mjsws = 0.29781 cjsws = {9.888891999999999E-11*sw_func_psd_nw_cj}
+ cjswgs = {2.39155046E-10*sw_func_psd_nw_cj} mjswgs = 0.9274 pbs = 0.6587
+ pbsws = 0.7418 pbswgs = 1.4338 xrcrg1 = 12
+ xrcrg2 = 1 rbpb = 50 rbpd = 50
+ rbps = 50 rbdb = 50 rbsb = 50
+ gbmin = 1E-12 tnom = 30 ute = 1.385810671525588
+ lute = -4.455758573125489E-6 wute = -6.101695540905441E-7 pute = 1.070097432373362E-12
+ kt1 = -0.639041164472424 lkt1 = 3.885591909686412E-7 wkt1 = 1.848465363671936E-7
+ pkt1 = -4.218824635666782E-13 kt1l = 0 kt2 = 0.054029277838872
+ lkt2 = -1.730179940720891E-7 wkt2 = -6.08197590947772E-8 pkt2 = 9.487868920509252E-14
+ ua1 = 7.897588967966098E-9 lua1 = -1.667562845925237E-14 wua1 = -3.819449800359685E-15
+ pua1 = 8.089209477761397E-21 ub1 = -6.528041614985322E-18 lub1 = 1.530911058287208E-23
+ wub1 = 3.671267371420774E-24 pub1 = -7.993205785764078E-30 uc1 = -3.281367055528903E-10
+ luc1 = 8.28879897592411E-16 wuc1 = 1.027620520043811E-16 puc1 = -2.458048002778201E-22
+ at = 1.248741640863949E5 lat = -0.316469148996462 wat = -0.020818996820791
+ pat = 1.194297209311976E-7 prt = 0 njs = 1.3632
+ xtis = 5.2 tpb = 2.0386E-3 tpbsw = 1.246E-3
+ tpbswg = 0 tcj = 1.2407E-3 tcjsw = 3.7357E-4
+ tcjswg = 2E-12 tvoff = 0 tvfbsdoff = 0
+ saref = 3E-6 sbref = 3E-6 wlod = 0
+ ku0 = 4.5E-8 kvsat = 0.5 kvth0 = 3.29E-8
+ tku0 = 0 llodku0 = 0 wlodku0 = 1
+ llodvth = 0 wlodvth = 1 lku0 = 0
+ wku0 = 2.5E-7 pku0 = 0 lkvth0 = 0
+ wkvth0 = 2E-7 pkvth0 = 0 stk2 = 0
+ lodk2 = 1 steta0 = 0 lodeta0 = 1

.model pshort_model.36 pmos
+ level = 54 lmin = 1E-6 lmax = 2E-6 wmin = 5.5E-7
+ wmax = 1E-6 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 4.23E-9
+ toxm = 4.23E-9 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 9.999999999999999E22 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {7.3039E-9+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {-1.3994E-8-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = -5.722E-9 dwb = -1.7864E-8 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = -0.97437499225458 lvth0 = -3.37450612343046E-8
+ wvth0 = -5.431924724776384E-8 pvth0 = 5.21896065766968E-14 k1 = 0.53590406200807
+ lk1 = -1.229448607405876E-7 wk1 = -6.585275404395844E-8 pk1 = 1.054838075947878E-13
+ k2 = -0.010300709913393 lk2 = 2.625822787125839E-8 wk2 = 1.435993576254715E-8
+ pk2 = -2.261320685988812E-14 k3 = -15.845 k3b = 2
+ w0 = 0 lpe0 = 0 lpeb = 0
+ vbm = -3 dvtp0 = 0 dvtp1 = 0
+ dvt0 = 4.4955 dvt1 = 0.294 dvt2 = 0.015
+ dvt0w = -4.9772 dvt1w = 1.1472E6 dvt2w = -8.96E-3
+ vfbsdoff = 0 u0 = -2.213911905194913E-3 lu0 = 1.50635077236042E-8
+ wu0 = 9.08205842231567E-9 pu0 = -1.317599277363353E-14 ua = -3.367067277808776E-9
+ lua = 3.781937036812744E-15 wua = 2.037873645442569E-15 pua = -3.187663906263714E-21
+ ub = 2.561415001513062E-18 lub = -2.316635270131664E-24 wub = -1.219882815046394E-24
+ pub = 1.921547836650994E-30 uc = 3.922729640764734E-11 luc = -1.192742692620113E-16
+ wuc = -7.933408768584968E-17 puc = 1.100391097082805E-22 ud = 0
+ up = 0 lp = 1 eu = 1.67
+ vsat = 2.004709379928953E5 lvsat = -0.247162471520137 wvsat = -0.119939300160125
+ pvsat = 1.92961168892021E-7 a0 = 2.155572234243662 la0 = -2.468249519082085E-6
+ wa0 = -5.648603575014886E-7 pa0 = 1.388004524694464E-12 ags = -1.644758902101962
+ lags = 3.918417068132512E-6 wags = 1.251652914407872E-6 pags = -2.230705964075328E-12
+ b0 = 1.323716012429543E-7 lb0 = -8.827069251476402E-14 wb0 = -1.304379433663175E-13
+ pb0 = 8.698125189264686E-20 b1 = -6.137833485215178E-10 lb1 = 6.923301483330344E-16
+ wb1 = 6.048173241229852E-16 pb1 = -6.82216727992215E-22 keta = 0.077328547773627
+ lketa = -1.654003674474182E-7 wketa = -4.748793651751838E-8 pketa = 9.513807518795559E-14
+ a1 = 0 a2 = 0.310776216094578 la2 = 9.921399630747894E-7
+ wa2 = 4.820773007148888E-7 pa2 = -9.776469809221857E-13 rdsw = 547.88
+ rdswmin = 0 rdw = 0 rdwmin = 0
+ rsw = 0 rswmin = 0 prwb = -0.32348
+ prwg = 0.1376 wr = 1 voff = -0.238478313326255
+ lvoff = 2.626694580201212E-8 wvoff = -8.053978557794696E-9 pvoff = -2.15162258443572E-14
+ voffl = 0 minv = 0 nfactor = 0.397978937900661
+ lnfactor = 1.748368703521905E-6 wnfactor = 1.086449076548965E-6 pnfactor = -1.399162165275983E-12
+ eta0 = 0.420229332503058 leta0 = -8.512060495642112E-7 weta0 = -4.941292332327609E-7
+ peta0 = 1.00208815544524E-12 etab = -0.187061479259446 letab = 3.783444345836008E-7
+ wetab = 1.904205373249662E-7 petab = -3.861705611059984E-13 dsub = -0.415314237929067
+ ldsub = 1.369529170749292E-6 wdsub = 3.615579755361666E-7 pdsub = -7.332352356916394E-13
+ cit = 1E-5 cdsc = 1.3E-4 cdscb = 7.8E-4
+ cdscd = 0 pclm = 0.832353444955653 lpclm = -8.490211770819548E-7
+ wpclm = -4.923899776324068E-7 ppclm = 8.758333822996524E-13 pdiblc1 = 0.40809150107188
+ lpdiblc1 = -3.668934707575991E-8 wpdiblc1 = -9.965887622218775E-9 ppdiblc1 = 2.021070050720821E-14
+ pdiblc2 = 2.996531676710831E-4 lpdiblc2 = -3.499802243770258E-10 wpdiblc2 = -8.341657112837738E-11
+ ppdiblc2 = 3.448677832553711E-16 pdiblcb = -1.157773472794311 lpdiblcb = 1.40908942870359E-6
+ wpdiblcb = 7.165534330797065E-7 ppdiblcb = -9.776469809221857E-13 drout = 0.170929482856047
+ ldrout = 7.890303399217308E-7 wdrout = 2.757802741494132E-8 pdrout = -5.592790866117202E-14
+ pscbe1 = 7.98527791097688E8 lpscbe1 = 2.985621987381887 wpscbe1 = 1.450703169108797
+ ppscbe1 = -2.94200861851461E-6 pscbe2 = 1.071579923042003E-8 lpscbe2 = -3.101498653131511E-15
+ wpscbe2 = -3.49280520629974E-16 ppscbe2 = 1.079397056932132E-21 pvag = 0
+ delta = 0.01 fprout = 0 pdits = 0
+ pditsl = 0 pditsd = 0 lambda = 0
+ vtl = 0 lc = 5E-9 xn = 3
+ alpha0 = -9.822235348678354E-11 lalpha0 = 2.037702007161716E-16 walpha0 = 1.583389808401636E-18
+ palpha0 = -1.627705722359182E-24 alpha1 = -1.02810558040378E-10 lalpha1 = 2.08486819938812E-16
+ walpha1 = 5.743345007077588E-21 palpha1 = -5.904089747135675E-27 beta0 = -4.260470984952272
+ lbeta0 = 1.472414803183139E-5 wbeta0 = 1.176840960019603E-6 pbeta0 = -2.386619344828234E-12
+ aigbacc = 0.43 bigbacc = 0.054 cigbacc = 0.075
+ nigbacc = 1 aigbinv = 0.35 bigbinv = 0.03
+ cigbinv = 6E-3 eigbinv = 1.1 nigbinv = 3
+ aigc = 0.43 bigc = 0.054 cigc = 0.075
+ aigsd = 0.43 bigsd = 0.054 cigsd = 0.075
+ dlcig = 0 nigc = 1 poxedge = 1
+ pigcd = 1 ntox = 1 toxref = 4.23E-9
+ agidl = 7.992204482993586E-10 lagidl = -1.366998070076286E-15 wagidl = -3.924842752884688E-16
+ pagidl = 1.042208074571915E-21 bgidl = 1E9 cgidl = 300
+ egidl = 0.1 noia = 1.5E42 noib = 0
+ noic = 0 em = 4.1E7 af = 1
+ ef = 1 kf = 0 lintnoi = -2E-7
+ tnoia = 2.5E7 tnoib = 0 ntnoi = 1
+ rnoia = 0.69 rnoib = 0.34 xpart = 0
+ cgso = {5.248925E-11/sw_func_tox_lv_ratio} cgdo = {5.248925E-11/sw_func_tox_lv_ratio} cgbo = {0/sw_func_tox_lv_ratio}
+ ckappas = 0.6 cf = 1.2E-11 clc = 1E-7
+ cle = 0.6 dlc = -3E-9 dwc = 0
+ vfbcv = -0.14469 noff = 3.9 voffcv = -0.10701
+ acde = 0.8 moin = 18.13 cgsl = {9.548271750000001E-12/sw_func_tox_lv_ratio}
+ cgdl = {9.548271750000001E-12/sw_func_tox_lv_ratio} ijthsrev = 0.1 ijthsfwd = 0.1
+ xjbvs = 1 bvs = 12.69 jss = 2.1483E-5
+ jsws = 8.040000000000001E-10 cjs = {sw_psd_nw_cj} mjs = 0.34629
+ mjsws = 0.29781 cjsws = {9.888891999999999E-11*sw_func_psd_nw_cj} cjswgs = {2.39155046E-10*sw_func_psd_nw_cj}
+ mjswgs = 0.9274 pbs = 0.6587 pbsws = 0.7418
+ pbswgs = 1.4338 xrcrg1 = 12 xrcrg2 = 1
+ rbpb = 50 rbpd = 50 rbps = 50
+ rbdb = 50 rbsb = 50 gbmin = 1E-12
+ tnom = 30 ute = 0.820533552469153 lute = -3.309383359004468E-6
+ wute = -1.388270738124446E-6 pute = 2.648077296379907E-12 kt1 = -0.385046571048059
+ lkt1 = -1.265387965608513E-7 wkt1 = -4.123537731923652E-8 pkt1 = 3.660894440643766E-14
+ kt1l = 0 kt2 = 7.298156265385096E-3 lkt2 = -7.824784029451676E-8
+ wkt2 = -3.34710799002653E-8 pkt2 = 3.941589598277275E-14 ua1 = 1.108865264176622E-9
+ lua1 = -2.908178252651758E-15 wua1 = -1.155454745078908E-15 pua1 = 2.686659473592642E-21
+ ub1 = 3.948956754725692E-19 lub1 = 1.269476833070958E-24 wub1 = 6.16885975125803E-25
+ pub1 = -1.798956966654634E-30 uc1 = 5.346529094308959E-11 luc1 = 5.499562792252179E-17
+ wuc1 = 2.289458638762197E-17 puc1 = -8.38345384166201E-23 at = -2.584541125061675E4
+ lat = -0.010811658847907 wat = 0.017126905172837 pat = 4.247588703894508E-8
+ prt = 0 njs = 1.3632 xtis = 5.2
+ tpb = 2.0386E-3 tpbsw = 1.246E-3 tpbswg = 0
+ tcj = 1.2407E-3 tcjsw = 3.7357E-4 tcjswg = 2E-12
+ tvoff = 0 tvfbsdoff = 0 saref = 3E-6
+ sbref = 3E-6 wlod = 0 ku0 = 4.5E-8
+ kvsat = 0.5 kvth0 = 3.29E-8 tku0 = 0
+ llodku0 = 0 wlodku0 = 1 llodvth = 0
+ wlodvth = 1 lku0 = 0 wku0 = 2.5E-7
+ pku0 = 0 lkvth0 = 0 wkvth0 = 2E-7
+ pkvth0 = 0 stk2 = 0 lodk2 = 1
+ steta0 = 0 lodeta0 = 1

.model pshort_model.37 pmos
+ level = 54 lmin = 5E-7 lmax = 1E-6 wmin = 5.5E-7
+ wmax = 1E-6 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 4.23E-9
+ toxm = 4.23E-9 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 9.999999999999999E22 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {7.3039E-9+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {-1.3994E-8-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = -5.722E-9 dwb = -1.7864E-8 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = -1.052142681599624 lvth0 = 4.619919020012746E-8
+ wvth0 = 7.917959881888625E-9 pvth0 = -1.178949550610038E-14 k1 = 0.352930576586212
+ lk1 = 6.51496865912579E-8 wk1 = 4.145470961424218E-8 pk1 = -4.826977356278529E-15
+ k2 = 0.028318272740247 lk2 = -1.344162286889093E-8 wk2 = -5.955573824548698E-9
+ pk2 = -1.729106790468637E-15 k3 = -15.845 k3b = 2
+ w0 = 0 lpe0 = 0 lpeb = 0
+ vbm = -3 dvtp0 = 0 dvtp1 = 0
+ dvt0 = 4.4955 dvt1 = 0.294 dvt2 = 0.015
+ dvt0w = -4.9772 dvt1w = 1.1472E6 dvt2w = -8.96E-3
+ vfbsdoff = 0 u0 = 0.015637388673433 lu0 = -3.287415055618568E-9
+ wu0 = -5.164717753982268E-9 pu0 = 1.469522174286634E-15 ua = 9.98771106986636E-10
+ lua = -7.060924326963218E-16 wua = -1.354888914038988E-15 pua = 3.000552917326114E-22
+ ub = -8.31197463605112E-20 lub = 4.019147162653941E-25 wub = 7.74365912286183E-25
+ pub = -1.285159240621666E-31 uc = -1.239392007187294E-10 luc = 4.845893178593849E-17
+ wuc = 4.618720362760979E-17 puc = -1.899527150646003E-23 ud = 0
+ up = 0 lp = 1 eu = 1.67
+ vsat = -1.772043013276464E5 lvsat = 0.141083142398508 wvsat = 0.139367155373281
+ pvsat = -7.360275571885395E-8 a0 = -1.742616559667892 la0 = 1.539041782793466E-6
+ wa0 = 1.653171692692884E-6 pa0 = -8.921058065207483E-13 ags = 2.46711240538198
+ lags = -3.085372935052897E-7 wags = -1.294843011735842E-6 pags = 3.870612900492961E-13
+ b0 = 9.901418678941586E-9 lb0 = 3.762718551885029E-14 wb0 = -9.756780735163353E-15
+ pb0 = -3.707753511822802E-20 b1 = 5.390810979638372E-10 lb1 = -4.928006682805528E-16
+ wb1 = -5.312063091010011E-16 pb1 = 4.856019346784442E-22 keta = -0.106238214481036
+ lketa = 2.330406134922794E-8 wketa = 6.273248935839687E-8 pketa = -1.816719996737477E-14
+ a1 = 0 a2 = 1.778447567810845 la2 = -5.166085744333121E-7
+ wa2 = -9.641546014297773E-7 pa2 = 5.090620596997052E-13 rdsw = 547.88
+ rdswmin = 0 rdw = 0 rdwmin = 0
+ rsw = 0 rswmin = 0 prwb = -0.32348
+ prwg = 0.1376 wr = 1 voff = -0.194013717710146
+ lvoff = -1.944212491620037E-8 wvoff = -4.704465572477757E-8 pvoff = 1.856572239517519E-14
+ voffl = 0 minv = 0 nfactor = 2.396422108663698
+ lnfactor = -3.060068947044488E-7 wnfactor = -6.495298862494808E-7 pnfactor = 3.854033767332661E-13
+ eta0 = -1.355858917006116 leta0 = 9.745913578722248E-7 weta0 = 9.882584664655217E-7
+ peta0 = -5.217886111921978E-13 etab = 0.372101557135284 letab = -1.964684568737441E-7
+ wetab = -3.80841067564762E-7 petab = 2.010795135813835E-13 dsub = 1.525156789700413
+ ldsub = -6.252517600014814E-7 wdsub = -6.986396470765472E-7 pdsub = 3.566351979827591E-13
+ cit = 1E-5 cdsc = 1.3E-4 cdscb = 7.8E-4
+ cdscd = 0 pclm = -0.642391681306558 lpclm = 6.669991157740828E-7
+ wpclm = 7.33774461116337E-7 ppclm = -3.846489467607912E-13 pdiblc1 = 0.653348915717859
+ lpdiblc1 = -2.888110262428502E-7 wpdiblc1 = -3.085306901286618E-8 ppdiblc1 = 4.168247233061705E-14
+ pdiblc2 = -1.379432587924257E-4 lpdiblc2 = 9.986365087034355E-11 wpdiblc2 = 1.773297554981966E-11
+ ppdiblc2 = 2.408872630647446E-16 pdiblcb = 0.212952088888889 wpdiblcb = -2.344761323648178E-7
+ drout = 0.666698216903657 ldrout = 2.793860305455967E-7 wdrout = 1.48636234100213E-7
+ pdrout = -1.803742924351511E-13 pscbe1 = 8.02944417804624E8 lpscbe1 = -1.554617267827806
+ wpscbe1 = -2.901406338217593 ppscbe1 = 1.53190772970283E-6 pscbe2 = -4.459582259469244E-9
+ lpscbe2 = 1.249861141389678E-14 wpscbe2 = 1.173736327090133E-14 ppscbe2 = -1.134552772103655E-20
+ pvag = 0 delta = 0.01 fprout = 0
+ pdits = 0 pditsl = 0 pditsd = 0
+ lambda = 0 vtl = 0 lc = 5E-9
+ xn = 3 alpha0 = 1E-10 alpha1 = 1E-10
+ beta0 = 11.185436212208492 lbeta0 = -1.15405921596351E-6 wbeta0 = -2.387204270820368E-6
+ pbeta0 = 1.277176383932486E-12 aigbacc = 0.43 bigbacc = 0.054
+ cigbacc = 0.075 nigbacc = 1 aigbinv = 0.35
+ bigbinv = 0.03 cigbinv = 6E-3 eigbinv = 1.1
+ nigbinv = 3 aigc = 0.43 bigc = 0.054
+ cigc = 0.075 aigsd = 0.43 bigsd = 0.054
+ cigsd = 0.075 dlcig = 0 nigc = 1
+ poxedge = 1 pigcd = 1 ntox = 1
+ toxref = 4.23E-9 agidl = -1.55307537140068E-9 lagidl = 1.051133805025518E-15
+ wagidl = 1.339274681192434E-15 pagidl = -7.380193515829752E-22 bgidl = 1E9
+ cgidl = 300 egidl = 0.1 noia = 1.5E42
+ noib = 0 noic = 0 em = 4.1E7
+ af = 1 ef = 1 kf = 0
+ lintnoi = -2E-7 tnoia = 2.5E7 tnoib = 0
+ ntnoi = 1 rnoia = 0.69 rnoib = 0.34
+ xpart = 0 cgso = {5.248925E-11/sw_func_tox_lv_ratio} cgdo = {5.248925E-11/sw_func_tox_lv_ratio}
+ cgbo = {0/sw_func_tox_lv_ratio} ckappas = 0.6 cf = 1.2E-11
+ clc = 1E-7 cle = 0.6 dlc = -3E-9
+ dwc = 0 vfbcv = -0.14469 noff = 3.9
+ voffcv = -0.10701 acde = 0.8 moin = 18.13
+ cgsl = {9.548271750000001E-12/sw_func_tox_lv_ratio} cgdl = {9.548271750000001E-12/sw_func_tox_lv_ratio} ijthsrev = 0.1
+ ijthsfwd = 0.1 xjbvs = 1 bvs = 12.69
+ jss = 2.1483E-5 jsws = 8.040000000000001E-10 cjs = {sw_psd_nw_cj}
+ mjs = 0.34629 mjsws = 0.29781 cjsws = {9.888891999999999E-11*sw_func_psd_nw_cj}
+ cjswgs = {2.39155046E-10*sw_func_psd_nw_cj} mjswgs = 0.9274 pbs = 0.6587
+ pbsws = 0.7418 pbswgs = 1.4338 xrcrg1 = 12
+ xrcrg2 = 1 rbpb = 50 rbpd = 50
+ rbps = 50 rbdb = 50 rbsb = 50
+ gbmin = 1E-12 tnom = 30 ute = -4.49096248907558
+ lute = 2.150770833751019E-6 wute = 2.257923225531147E-6 pute = -1.100166343930479E-12
+ kt1 = -0.508983522085384 lkt1 = 8.669018621064246E-10 wkt1 = -1.039733181517403E-8
+ pkt1 = 4.907803684807476E-15 kt1l = 0 kt2 = -0.108858432168539
+ lkt2 = 4.115973873649652E-8 wkt2 = 3.528623023832586E-8 pkt2 = -3.126579375197731E-14
+ ua1 = -4.430175614938374E-9 lua1 = 2.785889302587908E-15 wua1 = 3.299532786318834E-15
+ pua1 = -1.893014248833859E-21 ub1 = 2.674831976509397E-18 lub1 = -1.074270325159287E-24
+ wub1 = -2.237342598328365E-24 pub1 = 1.13515575611337E-30 uc1 = 1.942332745370531E-10
+ luc1 = -8.97121699962696E-17 wuc1 = -1.205983566903627E-16 puc1 = 6.367448515223122E-23
+ at = -1.422685803096367E5 lat = 0.108869961866737 wat = 0.119050074809943
+ pat = -6.229990826996469E-8 prt = 0 njs = 1.3632
+ xtis = 5.2 tpb = 2.0386E-3 tpbsw = 1.246E-3
+ tpbswg = 0 tcj = 1.2407E-3 tcjsw = 3.7357E-4
+ tcjswg = 2E-12 tvoff = 0 tvfbsdoff = 0
+ saref = 2.75E-6 sbref = 2.74E-6 wlod = 0
+ ku0 = 4.5E-8 kvsat = 0.5 kvth0 = 3.29E-8
+ tku0 = 0 llodku0 = 0 wlodku0 = 1
+ llodvth = 0 wlodvth = 1 lku0 = 0
+ wku0 = 2.5E-7 pku0 = 0 lkvth0 = 0
+ wkvth0 = 2E-7 pkvth0 = 0 stk2 = 0
+ lodk2 = 1 steta0 = 0 lodeta0 = 1

.model pshort_model.38 pmos
+ level = 54 lmin = 2.5E-7 lmax = 5E-7 wmin = 5.5E-7
+ wmax = 1E-6 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 4.23E-9
+ toxm = 4.23E-9 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 9.999999999999999E22 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {7.3039E-9+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {-1.3994E-8-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = -5.722E-9 dwb = -1.7864E-8 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = -1.0201764589423 lvth0 = 2.932140823173268E-8
+ wvth0 = 3.032009294931167E-8 pvth0 = -2.361755294010301E-14 k1 = 1.212301265021453
+ lk1 = -3.885877244542881E-7 wk1 = -7.708539083351195E-7 pk1 = 4.24062225217569E-13
+ k2 = -0.313455798341035 lk2 = 1.670109853731726E-7 wk2 = 3.189756309469768E-7
+ pk2 = -1.732888837353768E-13 k3 = -15.845 k3b = 2
+ w0 = 0 lpe0 = 0 lpeb = 0
+ vbm = -3 dvtp0 = 0 dvtp1 = 0
+ dvt0 = 4.4955 dvt1 = 0.294 dvt2 = 0.015
+ dvt0w = -4.9772 dvt1w = 1.1472E6 dvt2w = -8.96E-3
+ vfbsdoff = 0 u0 = 0.011258568707022 lu0 = -9.754506591932495E-10
+ wu0 = -1.969690631352895E-9 pu0 = -2.174138061362037E-16 ua = -1.757997990310847E-10
+ lua = -8.593308916983746E-17 wua = -4.425364651600804E-16 pua = -1.816558530460651E-22
+ ub = 8.506642254090864E-19 lub = -9.111201542129236E-26 wub = 3.832937378058431E-27
+ pub = 2.783162402936243E-31 uc = -6.784392879138671E-11 luc = 1.884130135156466E-17
+ wuc = 2.143042725988434E-17 puc = -5.923990665617403E-24 ud = 0
+ up = 0 lp = 1 eu = 1.67
+ vsat = -1.157551221391331E5 lvsat = 0.108638713177123 wvsat = 0.107919543353693
+ pvsat = -5.699879394385607E-8 a0 = 1.352455150621745 la0 = -9.511893937893853E-8
+ wa0 = 1.401391443712776E-7 pa0 = -9.324277739752009E-14 ags = 5.429764176989441
+ lags = -1.87278187709277E-6 wags = -3.080833087898378E-6 pags = 1.330042618382201E-12
+ b0 = 2.0706977201689E-7 lb0 = -6.647533902334643E-14 wb0 = -2.040449382012218E-13
+ pb0 = 6.55042805659612E-20 b1 = 2.50420392426451E-9 lb1 = -1.530361939093392E-15
+ wb1 = -2.467623014179638E-15 pb1 = 1.508006717959504E-21 keta = -0.139943697649754
+ lketa = 4.11001519965134E-8 wketa = 7.940456709413033E-8 pketa = -2.696985694690921E-14
+ a1 = 0 a2 = 1.472708584158838 la2 = -3.551820599328568E-7
+ wa2 = -3.601629288316858E-7 pa2 = 1.901617044679841E-13 rdsw = 547.88
+ rdswmin = 0 rdw = 0 rdwmin = 0
+ rsw = 0 rswmin = 0 prwb = -0.32348
+ prwg = 0.1376 wr = 1 voff = -0.300938880151905
+ lvoff = 3.701307775109888E-8 wvoff = 1.037604887137283E-7 pvoff = -6.105758420662265E-14
+ voffl = 0 minv = 0 nfactor = 3.117728783693762
+ lnfactor = -6.868481634402219E-7 wnfactor = -1.173022321772212E-6 pnfactor = 6.618011007800417E-13
+ eta0 = 0.079408144954019 leta0 = 2.167875723620175E-7 weta0 = 4.045940113458406E-7
+ peta0 = -2.136207828624677E-13 etab = -0.029371376551866 letab = 1.550443443786674E-8
+ wetab = 2.899780027777294E-8 petab = -1.531049057306078E-14 dsub = -0.465103663913313
+ ldsub = 4.255818763811225E-7 wdsub = 4.307839860384208E-7 pdsub = -2.396869272183466E-13
+ cit = 1E-5 cdsc = 1.3E-4 cdscb = 7.8E-4
+ cdscd = 0 pclm = 0.576833570663483 lpclm = 2.326281343692475E-8
+ wpclm = 3.669979530686447E-8 ppclm = -1.66018881093795E-14 pdiblc1 = -0.664867106707794
+ lpdiblc1 = 4.071912150056254E-7 wpdiblc1 = 4.718780866635611E-7 ppdiblc1 = -2.237535450926684E-13
+ pdiblc2 = -0.022031802514091 lpdiblc2 = 1.165955861135688E-8 wpdiblc2 = 1.069082705527065E-8
+ ppdiblc2 = -5.394378333898895E-15 pdiblcb = 0.898377265891201 lpdiblcb = -3.618962683550964E-7
+ wpdiblcb = -6.907469899516348E-7 ppdiblcb = 2.409055375555483E-13 drout = 2.797434955052282
+ ldrout = -8.456173983560197E-7 wdrout = -1.148464694588167E-6 pdrout = 5.044794327011693E-13
+ pscbe1 = 8E8 pscbe2 = 3.058951776577069E-8 lpscbe2 = -6.006892810229594E-15
+ wpscbe2 = -2.084385848787991E-14 ppscbe2 = 5.856966392938838E-21 pvag = 0
+ delta = 0.01 fprout = 0 pdits = 0
+ pditsl = 0 pditsd = 0 lambda = 0
+ vtl = 0 lc = 5E-9 xn = 3
+ alpha0 = 1E-10 alpha1 = 1E-10 beta0 = 6.645299395366361
+ lbeta0 = 1.243078541687334E-6 wbeta0 = 2.065436881187451E-6 pbeta0 = -1.073764712633819E-12
+ aigbacc = 0.43 bigbacc = 0.054 cigbacc = 0.075
+ nigbacc = 1 aigbinv = 0.35 bigbinv = 0.03
+ cigbinv = 6E-3 eigbinv = 1.1 nigbinv = 3
+ aigc = 0.43 bigc = 0.054 cigc = 0.075
+ aigsd = 0.43 bigsd = 0.054 cigsd = 0.075
+ dlcig = 0 nigc = 1 poxedge = 1
+ pigcd = 1 ntox = 1 toxref = 4.23E-9
+ agidl = 2.683373306853128E-9 lagidl = -1.185660259708353E-15 wagidl = -1.96633011466548E-15
+ pagidl = 1.007300313372453E-21 bgidl = 3.246615685604725E8 lbgidl = 356.57058773889327
+ wbgidl = 361.5709285529579 pbgidl = -1.909051114248191E-4 cgidl = 300
+ egidl = 0.1 noia = 1.5E42 noib = 0
+ noic = 0 em = 4.1E7 af = 1
+ ef = 1 kf = 0 lintnoi = -2E-7
+ tnoia = 2.5E7 tnoib = 0 ntnoi = 1
+ rnoia = 0.69 rnoib = 0.34 xpart = 0
+ cgso = {5.248925E-11/sw_func_tox_lv_ratio} cgdo = {5.248925E-11/sw_func_tox_lv_ratio} cgbo = {0/sw_func_tox_lv_ratio}
+ ckappas = 0.6 cf = 1.2E-11 clc = 1E-7
+ cle = 0.6 dlc = -3E-9 dwc = 0
+ vfbcv = -0.14469 noff = 3.9 voffcv = -0.10701
+ acde = 0.8 moin = 18.13 cgsl = {9.548271750000001E-12/sw_func_tox_lv_ratio}
+ cgdl = {9.548271750000001E-12/sw_func_tox_lv_ratio} ijthsrev = 0.1 ijthsfwd = 0.1
+ xjbvs = 1 bvs = 12.69 jss = 2.1483E-5
+ jsws = 8.040000000000001E-10 cjs = {sw_psd_nw_cj} mjs = 0.34629
+ mjsws = 0.29781 cjsws = {9.888891999999999E-11*sw_func_psd_nw_cj} cjswgs = {2.39155046E-10*sw_func_psd_nw_cj}
+ mjswgs = 0.9274 pbs = 0.6587 pbsws = 0.7418
+ pbswgs = 1.4338 xrcrg1 = 12 xrcrg2 = 1
+ rbpb = 50 rbpd = 50 rbps = 50
+ rbdb = 50 rbsb = 50 gbmin = 1E-12
+ tnom = 30 ute = -0.430498376869161 lute = 6.894508075377106E-9
+ wute = 1.26436376899013E-7 pute = 2.523313430510399E-14 kt1 = -0.674465132042276
+ lkt1 = 8.82392061400263E-8 wkt1 = 1.67535671141973E-7 pkt1 = -8.903868668053067E-14
+ kt1l = 0 kt2 = -0.18118469884309 lkt2 = 7.934713962545915E-8
+ wkt2 = 8.296189518424284E-8 pkt2 = -5.643797273544212E-14 ua1 = 1.00710868423836E-9
+ lua1 = -8.493155996581679E-17 wua1 = -2.759344709053845E-16 pua1 = -5.210442626558542E-24
+ ub1 = 7.760971200961845E-19 lub1 = -7.176110579138859E-26 wub1 = -9.802819617284754E-26
+ pub1 = 5.623423548082431E-33 uc1 = 8.254555810270692E-11 luc1 = -3.074239597153201E-17
+ wuc1 = -3.135449009881869E-17 puc1 = 1.655479451829508E-23 at = 5.055567808115046E4
+ lat = 7.061067327502334E-3 wat = 0.012528399217418 pat = -6.05774181721823E-9
+ prt = 0 njs = 1.3632 xtis = 5.2
+ tpb = 2.0386E-3 tpbsw = 1.246E-3 tpbswg = 0
+ tcj = 1.2407E-3 tcjsw = 3.7357E-4 tcjswg = 2E-12
+ tvoff = 0 tvfbsdoff = 0 saref = 1.75E-6
+ sbref = 1.74E-6 wlod = 0 ku0 = 4.5E-8
+ kvsat = 0.5 kvth0 = 3.29E-8 tku0 = 0
+ llodku0 = 0 wlodku0 = 1 llodvth = 0
+ wlodvth = 1 lku0 = 0 wku0 = 2.5E-7
+ pku0 = 0 lkvth0 = 0 wkvth0 = 2E-7
+ pkvth0 = 0 stk2 = 0 lodk2 = 1
+ steta0 = 0 lodeta0 = 1

.model pshort_model.39 pmos
+ level = 54 lmin = 1.8E-7 lmax = 2.5E-7 wmin = 5.5E-7
+ wmax = 1E-6 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 4.23E-9
+ toxm = 4.23E-9 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 9.999999999999999E22 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {7.3039E-9+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {-1.3994E-8-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = -5.722E-9 dwb = -1.7864E-8 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = -0.759152111552467 lvth0 = -4.324022805047237E-8
+ wvth0 = -1.379175063878794E-7 pvth0 = 2.315048082444412E-14 k1 = -3.75367803458284
+ lk1 = 9.918949290841099E-7 wk1 = 2.664959988195503E-6 pk1 = -5.310528082511856E-13
+ k2 = 1.610355053852367 lk2 = -3.677853458063667E-7 wk2 = -1.012730374903665E-6
+ pk2 = 1.969094054190315E-13 k3 = -15.845 k3b = 2
+ w0 = 0 lpe0 = 0 lpeb = 0
+ vbm = -3 dvtp0 = 0 dvtp1 = 0
+ dvt0 = 4.4955 dvt1 = 0.294 dvt2 = 0.015
+ dvt0w = -4.9772 dvt1w = 1.1472E6 dvt2w = -8.96E-3
+ vfbsdoff = 0 u0 = 0.020761959326326 lu0 = -3.61727921067228E-9
+ wu0 = -9.718503100784306E-9 pu0 = 1.936663074616096E-15 ua = 4.581535066979171E-9
+ lua = -1.408415093902296E-15 wua = -3.808546180268726E-15 pua = 7.540544556375571E-22
+ ub = -3.632311892981774E-18 lub = 1.155101549777946E-24 wub = 3.229686572256716E-24
+ pub = -6.18432359959024E-31 uc = -1.196736045753962E-12 luc = 3.141815345916997E-19
+ wuc = 7.252877480601724E-19 puc = -1.682103430044262E-25 ud = 0
+ up = 0 lp = 1 eu = 1.67
+ vsat = 7.598671453640368E5 lvsat = -0.134773769721548 wvsat = -0.356689069310772
+ pvsat = 7.215682507351317E-8 a0 = -0.778242254388763 la0 = 4.971893708451225E-7
+ wa0 = 7.622830271139354E-7 pa0 = -2.66191311073386E-13 ags = -6.695680835505494
+ lags = 1.497946331040672E-6 wags = 4.588675668019124E-6 pags = -8.019887816577936E-13
+ b0 = -3.206047469644445E-8 wb0 = 3.159214169417373E-14 b1 = -3.000932769022236E-9
+ wb1 = 2.957095743318907E-15 keta = -0.233431324503478 lketa = 6.708859041032622E-8
+ wketa = 1.115960684099219E-7 pketa = -3.591870801468346E-14 a1 = 0
+ a2 = -0.865925565527857 la2 = 2.949301700702484E-7 wa2 = 8.919235535642036E-7
+ pa2 = -1.579033126002844E-13 rdsw = 547.88 rdswmin = 0
+ rdw = 0 rdwmin = 0 rsw = 0
+ rswmin = 0 prwb = -0.32348 prwg = 0.1376
+ wr = 1 voff = 0.357565676486202 lvoff = -1.460432869396151E-7
+ wvoff = -3.97153294962022E-7 pvoff = 7.81904366898318E-14 voffl = 0
+ minv = 0 nfactor = -2.248780014860296 lnfactor = 8.049768844522235E-7
+ wnfactor = 2.758008679192087E-6 pnfactor = -4.309783451160218E-13 eta0 = 2.672118560677302
+ leta0 = -5.039548106840665E-7 weta0 = -1.334453205279314E-6 peta0 = 2.698134747927259E-13
+ etab = 0.231301797683951 letab = -5.695957992159956E-8 wetab = -1.357798353696715E-7
+ petab = 3.049571480530102E-14 dsub = 3.398440309066979 ldsub = -6.484369855797227E-7
+ wdsub = -1.68029646164005E-6 pdsub = 3.471681042708961E-13 cit = 1E-5
+ cdsc = 1.3E-4 cdscb = 7.8E-4 cdscd = 0
+ pclm = 0.758724971247986 lpclm = -2.730081322876008E-8 wpclm = -7.560192478793987E-8
+ ppclm = 1.461664245633496E-14 pdiblc1 = 2.814977781500222 lpdiblc1 = -5.601639057775447E-7
+ wpdiblc1 = -1.411875639999103E-6 ppdiblc1 = 2.999073858748324E-13 pdiblc2 = 0.076857963228805
+ lpdiblc2 = -1.583060958797938E-8 wpdiblc2 = -3.920328070674883E-8 ppdiblc2 = 8.475584894649376E-15
+ pdiblcb = -1.379415270921905 lpdiblcb = 2.713027233685052E-7 wpdiblcb = 6.983737616124749E-7
+ ppdiblcb = -1.452533619302554E-13 drout = -3.942172143870653 ldrout = 1.027912499859369E-6
+ wdrout = 2.646000416885626E-6 pdrout = -5.503363347072076E-13 pscbe1 = 8E8
+ pscbe2 = 7.818593645105025E-9 lpscbe2 = 3.231508442260115E-16 wpscbe2 = 8.476491828140012E-16
+ ppscbe2 = -1.730124414220216E-22 pvag = 0 delta = 0.01
+ fprout = 0 pdits = 0 pditsl = 0
+ pditsd = 0 lambda = 0 vtl = 0
+ lc = 5E-9 xn = 3 alpha0 = 1E-10
+ alpha1 = 1E-10 beta0 = 14.37531906463677 lbeta0 = -9.057741661338094E-7
+ wbeta0 = -3.541672548512263E-6 pbeta0 = 4.849444235095457E-13 aigbacc = 0.43
+ bigbacc = 0.054 cigbacc = 0.075 nigbacc = 1
+ aigbinv = 0.35 bigbinv = 0.03 cigbinv = 6E-3
+ eigbinv = 1.1 nigbinv = 3 aigc = 0.43
+ bigc = 0.054 cigc = 0.075 aigsd = 0.43
+ bigsd = 0.054 cigsd = 0.075 dlcig = 0
+ nigc = 1 poxedge = 1 pigcd = 1
+ ntox = 1 toxref = 4.23E-9 agidl = -1.581775763280667E-9
+ wagidl = 1.657208719285816E-15 bgidl = 3.392707140849234E9 lbgidl = -496.3092648105151
+ wbgidl = -1.281036740094982E3 pbgidl = 2.657201091672843E-4 cgidl = 300
+ egidl = 0.1 noia = 1.5E42 noib = 0
+ noic = 0 em = 4.1E7 af = 1
+ ef = 1 kf = 0 lintnoi = -2E-7
+ tnoia = 2.5E7 tnoib = 0 ntnoi = 1
+ rnoia = 0.69 rnoib = 0.34 xpart = 0
+ cgso = {5.248925E-11/sw_func_tox_lv_ratio} cgdo = {5.248925E-11/sw_func_tox_lv_ratio} cgbo = {0/sw_func_tox_lv_ratio}
+ ckappas = 0.6 cf = 1.2E-11 clc = 1E-7
+ cle = 0.6 dlc = -3E-9 dwc = 0
+ vfbcv = -0.14469 noff = 3.9 voffcv = -0.10701
+ acde = 0.8 moin = 18.13 cgsl = {9.548271750000001E-12/sw_func_tox_lv_ratio}
+ cgdl = {9.548271750000001E-12/sw_func_tox_lv_ratio} ijthsrev = 0.1 ijthsfwd = 0.1
+ xjbvs = 1 bvs = 12.69 jss = 2.1483E-5
+ jsws = 8.040000000000001E-10 cjs = {sw_psd_nw_cj} mjs = 0.34629
+ mjsws = 0.29781 cjsws = {9.888891999999999E-11*sw_func_psd_nw_cj} cjswgs = {2.39155046E-10*sw_func_psd_nw_cj}
+ mjswgs = 0.9274 pbs = 0.6587 pbsws = 0.7418
+ pbswgs = 1.4338 xrcrg1 = 12 xrcrg2 = 1
+ rbpb = 50 rbpd = 50 rbps = 50
+ rbdb = 50 rbsb = 50 gbmin = 1E-12
+ tnom = 30 ute = -0.20471603287926 lute = -5.58702741656875E-8
+ wute = 1.096033672184994E-7 pute = 2.991250900017059E-14 kt1 = 0.462819860899128
+ lkt1 = -2.279123744777688E-7 wkt1 = -5.917100310444782E-7 pkt1 = 1.220225075788765E-13
+ kt1l = 0 kt2 = 0.770550393763803 lkt2 = -1.852237952981458E-7
+ wkt2 = -4.767937345280687E-7 pkt2 = 9.916737525702397E-14 ua1 = 2.341444564514379E-9
+ lua1 = -4.558609226519869E-16 wua1 = -1.172645209855396E-15 pua1 = 2.440643822726771E-22
+ ub1 = 5.179525030933334E-19 wub1 = -7.779918071864657E-26 uc1 = -3.044427871710816E-11
+ luc1 = 6.67422786334744E-19 wuc1 = 2.948312689256572E-17 puc1 = -3.573329539058886E-25
+ at = 1.241812994444877E5 lat = -0.013405971904049 wat = -0.035082269617443
+ pat = 7.17745279084702E-9 prt = 0 njs = 1.3632
+ xtis = 5.2 tpb = 2.0386E-3 tpbsw = 1.246E-3
+ tpbswg = 0 tcj = 1.2407E-3 tcjsw = 3.7357E-4
+ tcjswg = 2E-12 tvoff = 0 tvfbsdoff = 0
+ saref = 1.04E-6 sbref = 1.04E-6 wlod = 0
+ ku0 = 4.5E-8 kvsat = 0.5 kvth0 = 3.29E-8
+ tku0 = 0 llodku0 = 0 wlodku0 = 1
+ llodvth = 0 wlodvth = 1 lku0 = 0
+ wku0 = 2.5E-7 pku0 = 0 lkvth0 = 0
+ wkvth0 = 2E-7 pkvth0 = 0 stk2 = 0
+ lodk2 = 1 steta0 = 0 lodeta0 = 1

.model pshort_model.40 pmos
+ level = 54 lmin = 1.5E-7 lmax = 1.8E-7 wmin = 5.5E-7
+ wmax = 1E-6 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 4.23E-9
+ toxm = 4.23E-9 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 9.999999999999999E22 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {7.3039E-9+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {-1.3994E-8-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = -5.722E-9 dwb = -1.7864E-8 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = -0.503869631600103 lvth0 = -9.633592049080457E-8
+ wvth0 = -2.745937549510313E-7 pvth0 = 5.157750041059694E-14 k1 = -3.775840560048527
+ lk1 = 9.965044684306671E-7 wk1 = 2.676825631462133E-6 pk1 = -5.335207196629255E-13
+ k2 = 1.704187750375173 lk2 = -3.87301420690752E-7 wk2 = -1.062967668726943E-6
+ pk2 = 2.073581596867473E-13 k3 = -15.845 k3b = 2
+ w0 = 0 lpe0 = 0 lpeb = 0
+ vbm = -3 dvtp0 = 0 dvtp1 = 0
+ dvt0 = 4.4955 dvt1 = 0.294 dvt2 = 0.015
+ dvt0w = -4.9772 dvt1w = 1.1472E6 dvt2w = -8.96E-3
+ vfbsdoff = 0 u0 = 8.798253837940365E-3 lu0 = -1.128972033553886E-9
+ wu0 = -3.313228499205336E-9 pu0 = 6.044428207828888E-16 ua = 6.420026475719322E-10
+ lua = -5.890396250546236E-16 wua = -1.699351251270962E-15 pua = 3.153672207451701E-22
+ ub = -9.89683774356381E-19 lub = 6.054666126412877E-25 wub = 1.814844090044007E-24
+ pub = -3.241621017685669E-31 uc = 2.758908759646666E-13 luc = 7.892806397285643E-21
+ wuc = -6.314521933799196E-20 puc = -4.225746981216834E-27 ud = 0
+ up = 0 lp = 1 eu = 1.67
+ vsat = 7.163505242805808E5 lvsat = -0.125722834735643 wvsat = -0.333390609812334
+ pvsat = 6.731102507935207E-8 a0 = 6.302834983750357 la0 = -9.75589721760957E-7
+ wa0 = -3.028870493783293E-6 pa0 = 5.223231274309867E-13 ags = 0.506399722222222
+ wags = 7.327379136400557E-7 b0 = -3.206047469644445E-8 wb0 = 3.159214169417373E-14
+ b1 = -3.000932769022191E-9 wb1 = 2.957095743318883E-15 keta = 0.446394902742544
+ lketa = -7.430710694211927E-8 wketa = -2.523775910130255E-7 pketa = 3.978344546137652E-14
+ a1 = 0 a2 = -3.510589910297408 la2 = 8.449886178101778E-7
+ wa2 = 2.307856215371932E-6 pa2 = -4.524003150643503E-13 rdsw = 547.88
+ rdswmin = 0 rdw = 0 rdwmin = 0
+ rsw = 0 rswmin = 0 prwb = -0.32348
+ prwg = 0.1376 wr = 1 voff = -0.088298823512793
+ lvoff = -5.330882131382419E-8 wvoff = -1.584409194056601E-7 pvoff = 2.854112712261522E-14
+ voffl = 0 minv = 0 nfactor = -3.805616460735225
+ lnfactor = 1.128780183156858E-6 wnfactor = 3.591526768989246E-6 pnfactor = -6.043401055767535E-13
+ eta0 = -1.451959625358182 leta0 = 3.538039630730817E-7 weta0 = 8.73546087714233E-7
+ peta0 = -1.89423882158416E-13 etab = -0.452508249858103 letab = 8.526470424657713E-8
+ wetab = 2.303267303659732E-7 petab = -4.565005758892427E-14 dsub = 0.32233240511297
+ ldsub = -8.64345485213643E-9 wdsub = -3.337228350472418E-8 pdsub = 4.627638308885999E-15
+ cit = 1E-5 cdsc = 1.3E-4 cdscb = 7.8E-4
+ cdscd = 0 pclm = 2.814153489590923 lpclm = -4.548052799018708E-7
+ wpclm = -1.176062321166305E-6 ppclm = 2.434991993782784E-13 pdiblc1 = 1.846277151208034
+ lpdiblc1 = -3.586857990843329E-7 wpdiblc1 = -8.932408784055816E-7 ppdiblc1 = 1.92037579080519E-13
+ pdiblc2 = 0.025232687084711 lpdiblc2 = -5.093171653321575E-9 wpdiblc2 = -1.156351053635486E-8
+ ppdiblc2 = 2.726844376449476E-15 pdiblcb = -1.049060524715446 lpdiblcb = 2.025929004145163E-7
+ wpdiblcb = 5.215044072605574E-7 ppdiblcb = -1.084666586573088E-13 drout = 1
+ pscbe1 = 8E8 pscbe2 = 9.530843849774069E-9 lpscbe2 = -3.297665134269347E-17
+ wpscbe2 = -6.90762212142083E-17 ppscbe2 = 1.765544191099761E-23 pvag = 0
+ delta = 0.01 fprout = 0 pdits = 0
+ pditsl = 0 pditsd = 0 lambda = 0
+ vtl = 0 lc = 5E-9 xn = 3
+ alpha0 = 1E-10 alpha1 = 1E-10 beta0 = 30.04242357294406
+ lbeta0 = -4.164343898607627E-6 wbeta0 = -1.192971809884482E-5 pbeta0 = 2.229557241432114E-12
+ aigbacc = 0.43 bigbacc = 0.054 cigbacc = 0.075
+ nigbacc = 1 aigbinv = 0.35 bigbinv = 0.03
+ cigbinv = 6E-3 eigbinv = 1.1 nigbinv = 3
+ aigc = 0.43 bigc = 0.054 cigc = 0.075
+ aigsd = 0.43 bigsd = 0.054 cigsd = 0.075
+ dlcig = 0 nigc = 1 poxedge = 1
+ pigcd = 1 ntox = 1 toxref = 4.23E-9
+ agidl = -1.223357045933443E-8 lagidl = 2.215445475242831E-15 wagidl = 7.360096515554372E-15
+ pagidl = -1.186132226970305E-21 bgidl = 1.044836933347849E9 lbgidl = -7.9804360927169
+ wbgidl = -24.0053443863581 pbgidl = 4.272663236639106E-6 cgidl = 300
+ egidl = 0.1 noia = 1.5E42 noib = 0
+ noic = 0 em = 4.1E7 af = 1
+ ef = 1 kf = 0 lintnoi = -2E-7
+ tnoia = 2.5E7 tnoib = 0 ntnoi = 1
+ rnoia = 0.69 rnoib = 0.34 xpart = 0
+ cgso = {5.248925E-11/sw_func_tox_lv_ratio} cgdo = {5.248925E-11/sw_func_tox_lv_ratio} cgbo = {0/sw_func_tox_lv_ratio}
+ ckappas = 0.6 cf = 1.2E-11 clc = 1E-7
+ cle = 0.6 dlc = -3E-9 dwc = 0
+ vfbcv = -0.14469 noff = 3.9 voffcv = -0.10701
+ acde = 0.8 moin = 18.13 cgsl = {9.548271750000001E-12/sw_func_tox_lv_ratio}
+ cgdl = {9.548271750000001E-12/sw_func_tox_lv_ratio} ijthsrev = 0.1 ijthsfwd = 0.1
+ xjbvs = 1 bvs = 12.69 jss = 2.1483E-5
+ jsws = 8.040000000000001E-10 cjs = {sw_psd_nw_cj} mjs = 0.34629
+ mjsws = 0.29781 cjsws = {9.888891999999999E-11*sw_func_psd_nw_cj} cjswgs = {2.39155046E-10*sw_func_psd_nw_cj}
+ mjswgs = 0.9274 pbs = 0.6587 pbsws = 0.7418
+ pbswgs = 1.4338 xrcrg1 = 12 xrcrg2 = 1
+ rbpb = 50 rbpd = 50 rbps = 50
+ rbdb = 50 rbsb = 50 gbmin = 1E-12
+ tnom = 30 ute = -0.521797668864676 lute = 1.007890113964716E-8
+ wute = 2.793664018883304E-7 pute = -5.396165054738198E-15 kt1 = 0.298269324198017
+ lkt1 = -1.936878374503783E-7 wkt1 = -5.036109571888898E-7 pkt1 = 1.036989574058004E-13
+ kt1l = 0 kt2 = -0.12 ua1 = 7.06763278478338E-10
+ lua1 = -1.158668313319227E-16 wua1 = -2.9744959982573E-16 pua1 = 6.203419773382705E-23
+ ub1 = 1.428540947639438E-18 lub1 = -1.893914694042554E-25 wub1 = -5.653211313387639E-25
+ pub1 = 1.01398715465577E-31 uc1 = -1.184325362783377E-10 luc1 = 1.896792449997975E-17
+ wuc1 = 7.659135368243902E-17 puc1 = -1.015527882747806E-23 at = 5.53865206301635E5
+ lat = -0.102775068323453 wat = -0.265131681814286 pat = 5.502496993484404E-8
+ prt = 0 njs = 1.3632 xtis = 5.2
+ tpb = 2.0386E-3 tpbsw = 1.246E-3 tpbswg = 0
+ tcj = 1.2407E-3 tcjsw = 3.7357E-4 tcjswg = 2E-12
+ tvoff = 0 tvfbsdoff = 0 saref = 1.04E-6
+ sbref = 1.04E-6 wlod = 0 ku0 = 4.5E-8
+ kvsat = 0.5 kvth0 = 3.29E-8 tku0 = 0
+ llodku0 = 0 wlodku0 = 1 llodvth = 0
+ wlodvth = 1 lku0 = 0 wku0 = 2.5E-7
+ pku0 = 0 lkvth0 = 0 wkvth0 = 2E-7
+ pkvth0 = 0 stk2 = 0 lodk2 = 1
+ steta0 = 0 lodeta0 = 1

.model pshort_model.41 pmos
+ level = 54 lmin = 8E-6 lmax = 2.02E-5 wmin = 4.2E-7
+ wmax = 5.5E-7 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 4.23E-9
+ toxm = 4.23E-9 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 9.999999999999999E22 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {7.3039E-9+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {-1.3994E-8-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = -5.722E-9 dwb = -1.7864E-8 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = -1.138687303252638 lvth0 = 5.092372287315432E-7
+ wvth0 = 5.1804229778117E-8 pvth0 = -2.726416402124841E-13 k1 = 0.564852267623845
+ lk1 = -4.296987340294455E-7 wk1 = -4.614348220252891E-8 pk1 = 2.300573505492397E-13
+ k2 = -0.107540793365244 lk2 = 4.458514875610562E-7 wk2 = 5.642644497116667E-8
+ pk2 = -2.387054087985866E-13 k3 = -15.845 k3b = 2
+ w0 = 0 lpe0 = 0 lpeb = 0
+ vbm = -3 dvtp0 = 0 dvtp1 = 0
+ dvt0 = 4.4955 dvt1 = 0.294 dvt2 = 0.015
+ dvt0w = -4.9772 dvt1w = 1.1472E6 dvt2w = -8.96E-3
+ vfbsdoff = 0 u0 = 0.012464721800426 lu0 = -1.064874384839536E-8
+ wu0 = -2.142242591311882E-9 pu0 = 5.701254396228858E-15 ua = -1.439855629678346E-9
+ lua = 1.018915263249457E-15 wua = 2.814093358189571E-16 pua = -5.45519284404706E-22
+ ub = 2.551715618346924E-18 lub = -1.724085023379612E-24 wub = -8.204612245509899E-25
+ pub = 9.23061673654262E-31 uc = -3.941166329732871E-12 luc = -1.91850335556514E-16
+ wuc = -3.430171395445279E-17 puc = 1.027151732243402E-22 ud = 0
+ up = 0 lp = 1 eu = 1.67
+ vsat = -2.92319756188324E5 lvsat = 1.619137313240068 wvsat = 0.169618018447174
+ pvsat = -8.668734882376892E-7 a0 = -0.504927130230126 la0 = 1.368554892140962E-5
+ wa0 = 9.40073175545554E-7 pa0 = -7.327136145241125E-12 ags = 0.729584329189763
+ lags = -3.726808607140947E-6 wags = -2.648163801861434E-7 pags = 1.995304259156127E-12
+ b0 = 1.489331376709344E-7 lb0 = -4.589059822613021E-12 wb0 = -1.200076999457444E-13
+ pb0 = 2.456946834360395E-18 b1 = -2.755327509253987E-9 lb1 = -6.268216499639497E-14
+ wb1 = 1.468247527910013E-15 pb1 = 3.35595422181829E-20 keta = -0.077079581257084
+ lketa = 6.123879136515651E-7 wketa = 4.523378095030386E-8 pketa = -3.278677123433215E-13
+ a1 = 0 a2 = -0.238319505333507 la2 = 8.335616528983335E-6
+ wa2 = 5.559081642634184E-7 pa2 = -4.462824071808752E-12 rdsw = 547.88
+ rdswmin = 0 rdw = 0 rdwmin = 0
+ rsw = 0 rswmin = 0 prwb = -0.32348
+ prwg = 0.1376 wr = 1 voff = -0.398443040851589
+ lvoff = -3.408431509574341E-7 wvoff = 5.902676564120999E-8 pvoff = 1.824847644460328E-13
+ voffl = 0 minv = 0 nfactor = 4.408182466368965
+ lnfactor = -2.702919550449833E-5 wnfactor = -1.473804501211166E-6 pnfactor = 1.447122044538347E-11
+ eta0 = 0.08 etab = -0.07 dsub = 0.56
+ cit = -4.310375541461448E-7 lcit = 2.089126949619884E-10 wcit = 5.584696144396923E-12
+ pcit = -1.118502273636279E-16 cdsc = 1.3E-4 cdscb = 7.8E-4
+ cdscd = 0 pclm = 1.285152216388717 lpclm = -2.560425569186176E-5
+ wpclm = -6.871287645432993E-7 ppclm = 1.370831878422839E-11 pdiblc1 = 0.39
+ pdiblc2 = -8.08025555849982E-3 lpdiblc2 = 8.008727868616044E-8 wpdiblc2 = 4.774697555664214E-9
+ ppdiblc2 = -4.287810432779655E-14 pdiblcb = -0.225 drout = 0.56
+ pscbe1 = 1.539133660722752E9 lpscbe1 = -5.949229377003598E3 wpscbe1 = -401.0282196934259
+ ppscbe1 = 3.185171004458586E-3 pscbe2 = 7.465748917323658E-9 lpscbe2 = 1.727222892057942E-14
+ wpscbe2 = 1.098661994882948E-15 ppscbe2 = -9.247416640692642E-21 pvag = 0
+ delta = 0.01 fprout = 0 pdits = 0
+ pditsl = 0 pditsd = 0 lambda = 0
+ vtl = 0 lc = 5E-9 xn = 3
+ alpha0 = 6.204609049290764E-10 lalpha0 = -4.178253899239767E-15 walpha0 = -2.786507089039691E-16
+ palpha0 = 2.237004547272557E-21 alpha1 = 6.204609049290764E-10 lalpha1 = -4.178253899239767E-15
+ walpha1 = -2.786507089039691E-16 palpha1 = 2.237004547272557E-21 beta0 = -133.7157207852456
+ lbeta0 = 1.051847483328041E-3 wbeta0 = 7.319653052579836E-5 pbeta0 = -5.631509381634632E-10
+ aigbacc = 0.43 bigbacc = 0.054 cigbacc = 0.075
+ nigbacc = 1 aigbinv = 0.35 bigbinv = 0.03
+ cigbinv = 6E-3 eigbinv = 1.1 nigbinv = 3
+ aigc = 0.43 bigc = 0.054 cigc = 0.075
+ aigsd = 0.43 bigsd = 0.054 cigsd = 0.075
+ dlcig = 0 nigc = 1 poxedge = 1
+ pigcd = 1 ntox = 1 toxref = 4.23E-9
+ agidl = 3.658223308128976E-9 lagidl = -1.171946862434461E-14 wagidl = -1.33047965685461E-15
+ pagidl = 6.274512089618836E-21 bgidl = 1E9 cgidl = 300
+ egidl = 0.1 noia = 1.5E42 noib = 0
+ noic = 0 em = 4.1E7 af = 1
+ ef = 1 kf = 0 lintnoi = -2E-7
+ tnoia = 2.5E7 tnoib = 0 ntnoi = 1
+ rnoia = 0.69 rnoib = 0.34 xpart = 0
+ cgso = {5.248925E-11/sw_func_tox_lv_ratio} cgdo = {5.248925E-11/sw_func_tox_lv_ratio} cgbo = {0/sw_func_tox_lv_ratio}
+ ckappas = 0.6 cf = 1.2E-11 clc = 1E-7
+ cle = 0.6 dlc = -3E-9 dwc = 0
+ vfbcv = -0.14469 noff = 3.9 voffcv = -0.10701
+ acde = 0.8 moin = 18.13 cgsl = {9.548271750000001E-12/sw_func_tox_lv_ratio}
+ cgdl = {9.548271750000001E-12/sw_func_tox_lv_ratio} ijthsrev = 0.1 ijthsfwd = 0.1
+ xjbvs = 1 bvs = 12.69 jss = 2.1483E-5
+ jsws = 8.040000000000001E-10 cjs = {sw_psd_nw_cj} mjs = 0.34629
+ mjsws = 0.29781 cjsws = {9.888891999999999E-11*sw_func_psd_nw_cj} cjswgs = {2.39155046E-10*sw_func_psd_nw_cj}
+ mjswgs = 0.9274 pbs = 0.6587 pbsws = 0.7418
+ pbswgs = 1.4338 xrcrg1 = 12 xrcrg2 = 1
+ rbpb = 50 rbpd = 50 rbps = 50
+ rbdb = 50 rbsb = 50 gbmin = 1E-12
+ tnom = 30 ute = -4.249298659015382 wute = 1.600714881607296E-6
+ kt1 = -1.21334211937223 lkt1 = 2.089126949619883E-6 wkt1 = 3.68206412401361E-7
+ pkt1 = -1.118502273636278E-12 kt1l = 0 kt2 = -0.032318659992242
+ wkt2 = -1.07963657505018E-8 ua1 = -2.986271449305121E-9 wua1 = 1.461739268230657E-15
+ ub1 = 1.271706424121261E-18 wub1 = -4.16195920016415E-25 uc1 = -1.961641283609832E-10
+ luc1 = 2.841212651483038E-16 wuc1 = 1.094123368624892E-16 puc1 = -1.521163092145337E-22
+ at = -2.239974452424998E5 wat = 0.125280407002762 prt = 0
+ njs = 1.3632 xtis = 5.2 tpb = 2.0386E-3
+ tpbsw = 1.246E-3 tpbswg = 0 tcj = 1.2407E-3
+ tcjsw = 3.7357E-4 tcjswg = 2E-12 tvoff = 0
+ tvfbsdoff = 0 saref = 3E-6 sbref = 3E-6
+ wlod = 0 ku0 = 4.5E-8 kvsat = 0.5
+ kvth0 = 3.29E-8 tku0 = 0 llodku0 = 0
+ wlodku0 = 1 llodvth = 0 wlodvth = 1
+ lku0 = 0 wku0 = 2.5E-7 pku0 = 0
+ lkvth0 = 0 wkvth0 = 2E-7 pkvth0 = 0
+ stk2 = 0 lodk2 = 1 steta0 = 0
+ lodeta0 = 1

.model pshort_model.42 pmos
+ level = 54 lmin = 4E-6 lmax = 8E-6 wmin = 4.2E-7
+ wmax = 5.5E-7 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 4.23E-9
+ toxm = 4.23E-9 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 9.999999999999999E22 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {7.3039E-9+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {-1.3994E-8-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = -5.722E-9 dwb = -1.7864E-8 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = -1.234551487586235 lvth0 = 1.278833750191446E-6
+ wvth0 = 8.415936820877597E-8 pvth0 = -5.323883032721531E-13 k1 = 0.578837878854054
+ lk1 = -5.41975053158236E-7 wk1 = -4.485487895545063E-8 pk1 = 2.197124591449342E-13
+ k2 = -0.132263169415061 lk2 = 6.443224258204721E-7 wk2 = 6.060276907118605E-8
+ pk2 = -2.72232888557653E-13 k3 = -15.845 k3b = 2
+ w0 = 0 lpe0 = 0 lpeb = 0
+ vbm = -3 dvtp0 = 0 dvtp1 = 0
+ dvt0 = 4.4955 dvt1 = 0.294 dvt2 = 0.015
+ dvt0w = -4.9772 dvt1w = 1.1472E6 dvt2w = -8.96E-3
+ vfbsdoff = 0 u0 = 0.017775417652256 lu0 = -5.32829464185349E-8
+ wu0 = -4.183769062313019E-9 pu0 = 2.209060440710833E-14 ua = -1.582920818044586E-9
+ lua = 2.167440878671372E-15 wua = 3.219835807685366E-16 pua = -8.712488359689911E-22
+ ub = 4.070004504558712E-18 lub = -1.391288998242122E-23 wub = -1.40805029531154E-24
+ pub = 5.640219682651111E-30 uc = -8.460092785689411E-12 luc = -1.555724481952124E-16
+ wuc = -2.936307725107244E-17 puc = 6.306785703324319E-23 ud = 0
+ up = 0 lp = 1 eu = 1.67
+ vsat = -2.840682049354304E5 lvsat = 1.552893958800454 wvsat = 0.148225981579132
+ pvsat = -6.951384729654891E-7 a0 = 1.212122214148439 la0 = -9.890261066937046E-8
+ wa0 = 2.237991390065297E-8 pa0 = 4.009434692499956E-14 ags = 0.269181293730407
+ lags = -3.069856330966551E-8 wags = -1.782307363920002E-8 pags = 1.244495811694458E-14
+ b0 = -9.810130056321403E-7 lb0 = 4.48213425647034E-12 wb0 = 4.352869146828305E-13
+ pb0 = -2.000951668342428E-18 b1 = -2.129308866500654E-8 lb1 = 8.613875910885261E-14
+ wb1 = 1.130356694173345E-14 pb1 = -4.539828401215872E-20 keta = -0.014200424831381
+ lketa = 1.075948004158941E-7 wketa = 9.826451057164839E-9 pketa = -4.361809284916022E-14
+ a1 = 0 a2 = 0.8 rdsw = 547.88
+ rdswmin = 0 rdw = 0 rdwmin = 0
+ rsw = 0 rswmin = 0 prwb = -0.32348
+ prwg = 0.1376 wr = 1 voff = -0.711656369270886
+ lvoff = 2.173629691032743E-6 wvoff = 1.942318527494387E-7 pvoff = -9.029400523977819E-13
+ voffl = 0 minv = 0 nfactor = 0.010906908419421
+ lnfactor = 8.27207990741391E-6 wnfactor = 7.32772971930665E-7 pnfactor = -3.243157030069468E-12
+ eta0 = 0.08 etab = -0.07 dsub = 0.56
+ cit = 2.559200769230768E-5 wcit = -8.347839300801534E-12 cdsc = 1.3E-4
+ cdscb = 7.8E-4 cdscd = 0 pclm = -3.555185432400447
+ lpclm = 1.325391686856586E-5 wpclm = 1.68972497542161E-6 ppclm = -5.373034517965022E-12
+ pdiblc1 = 0.39 pdiblc2 = 3.587299874321525E-3 lpdiblc2 = -1.357971631786413E-8
+ wpdiblc2 = -1.252119549851064E-9 ppdiblc2 = 5.505111073474838E-15 pdiblcb = -0.225
+ drout = 0.56 pscbe1 = 7.570039765933372E8 lpscbe1 = 329.6983416311361
+ wpscbe1 = 12.378992737482543 ppscbe1 = -1.336571360501978E-4 pscbe2 = 9.362121947538264E-9
+ lpscbe2 = 2.048168990492944E-15 wpscbe2 = 5.019195386333884E-17 ppscbe2 = -8.303117330277136E-22
+ pvag = 0 delta = 0.01 fprout = 0
+ pdits = 0 pditsl = 0 pditsd = 0
+ lambda = 0 vtl = 0 lc = 5E-9
+ xn = 3 alpha0 = 4.264596194826362E-10 lalpha0 = -2.620813907691169E-15
+ walpha0 = -1.323441833532287E-16 palpha0 = 1.06245751582952E-21 alpha1 = 5.147216599585812E-10
+ lalpha1 = -3.329380509487571E-15 walpha1 = -1.681249261182612E-16 palpha1 = 1.349704889378287E-21
+ beta0 = -88.39895690002426 lbeta0 = 6.88045046658651E-4 wbeta0 = 3.779253602563093E-5
+ pbeta0 = -2.789280951640532E-10 aigbacc = 0.43 bigbacc = 0.054
+ cigbacc = 0.075 nigbacc = 1 aigbinv = 0.35
+ bigbinv = 0.03 cigbinv = 6E-3 eigbinv = 1.1
+ nigbinv = 3 aigc = 0.43 bigc = 0.054
+ cigc = 0.075 aigsd = 0.43 bigsd = 0.054
+ cigsd = 0.075 dlcig = 0 nigc = 1
+ poxedge = 1 pigcd = 1 ntox = 1
+ toxref = 4.23E-9 agidl = 6.649055255099138E-9 lagidl = -3.57298316046377E-14
+ wagidl = -2.353162170856222E-15 pagidl = 1.448459503983361E-20 bgidl = -3.338776031328201E8
+ lbgidl = 1.070835339141904E4 wbgidl = 540.7435760647408 pbgidl = -4.341082939724825E-3
+ cgidl = 300 egidl = 0.1 noia = 1.5E42
+ noib = 0 noic = 0 em = 4.1E7
+ af = 1 ef = 1 kf = 0
+ lintnoi = -2E-7 tnoia = 2.5E7 tnoib = 0
+ ntnoi = 1 rnoia = 0.69 rnoib = 0.34
+ xpart = 0 cgso = {5.248925E-11/sw_func_tox_lv_ratio} cgdo = {5.248925E-11/sw_func_tox_lv_ratio}
+ cgbo = {0/sw_func_tox_lv_ratio} ckappas = 0.6 cf = 1.2E-11
+ clc = 1E-7 cle = 0.6 dlc = -3E-9
+ dwc = 0 vfbcv = -0.14469 noff = 3.9
+ voffcv = -0.10701 acde = 0.8 moin = 18.13
+ cgsl = {9.548271750000001E-12/sw_func_tox_lv_ratio} cgdl = {9.548271750000001E-12/sw_func_tox_lv_ratio} ijthsrev = 0.1
+ ijthsfwd = 0.1 xjbvs = 1 bvs = 12.69
+ jss = 2.1483E-5 jsws = 8.040000000000001E-10 cjs = {sw_psd_nw_cj}
+ mjs = 0.34629 mjsws = 0.29781 cjsws = {9.888891999999999E-11*sw_func_psd_nw_cj}
+ cjswgs = {2.39155046E-10*sw_func_psd_nw_cj} mjswgs = 0.9274 pbs = 0.6587
+ pbsws = 0.7418 pbswgs = 1.4338 xrcrg1 = 12
+ xrcrg2 = 1 rbpb = 50 rbpd = 50
+ rbps = 50 rbdb = 50 rbsb = 50
+ gbmin = 1E-12 tnom = 30 ute = -9.063899478412027
+ lute = 3.865155760290643E-5 wute = 3.695535352900431E-6 pute = -1.681719360569563E-11
+ kt1 = -1.557516990827226 lkt1 = 4.85215868756213E-6 wkt1 = 4.809528619329921E-7
+ pkt1 = -2.023629417518819E-12 kt1l = 0 kt2 = 4.240563304569088E-3
+ lkt2 = -2.934970059161165E-7 wkt2 = -2.71115166916116E-8 pkt2 = 1.309778359734181E-13
+ ua1 = -7.637194127103772E-9 lua1 = 3.733755144629543E-14 wua1 = 3.611740093878616E-15
+ pua1 = -1.72601808282919E-20 ub1 = 3.057346988150791E-18 lub1 = -1.43351010203423E-23
+ wub1 = -1.333927170234678E-24 pub1 = 7.36753546397721E-30 uc1 = -9.265492982426406E-13
+ luc1 = -1.283243676716429E-15 wuc1 = 3.323919496946278E-17 puc1 = 4.594007598249798E-22
+ at = -5.097064152200856E5 lat = 2.293668182472419 wat = 0.249779710540662
+ pat = -9.994789148106225E-7 prt = 0 njs = 1.3632
+ xtis = 5.2 tpb = 2.0386E-3 tpbsw = 1.246E-3
+ tpbswg = 0 tcj = 1.2407E-3 tcjsw = 3.7357E-4
+ tcjswg = 2E-12 tvoff = 0 tvfbsdoff = 0
+ saref = 3E-6 sbref = 3E-6 wlod = 0
+ ku0 = 4.5E-8 kvsat = 0.5 kvth0 = 3.29E-8
+ tku0 = 0 llodku0 = 0 wlodku0 = 1
+ llodvth = 0 wlodvth = 1 lku0 = 0
+ wku0 = 2.5E-7 pku0 = 0 lkvth0 = 0
+ wkvth0 = 2E-7 pkvth0 = 0 stk2 = 0
+ lodk2 = 1 steta0 = 0 lodeta0 = 1

.model pshort_model.43 pmos
+ level = 54 lmin = 2E-6 lmax = 4E-6 wmin = 4.2E-7
+ wmax = 5.5E-7 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 4.23E-9
+ toxm = 4.23E-9 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 9.999999999999999E22 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {7.3039E-9+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {-1.3994E-8-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = -5.722E-9 dwb = -1.7864E-8 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = -0.764847969952619 lvth0 = -6.131263823945454E-7
+ wvth0 = -1.09062253378943E-7 pvth0 = 2.4590606982372E-13 k1 = 0.427985192937785
+ lk1 = 6.56577554802654E-8 wk1 = 2.545187203444779E-8 pk1 = -6.348229016136476E-14
+ k2 = 0.080197933921393 lk2 = -2.114683488855232E-7 wk2 = -3.182528466548735E-8
+ pk2 = 1.000662027570226E-13 k3 = -15.845 k3b = 2
+ w0 = 0 lpe0 = 0 lpeb = 0
+ vbm = -3 dvtp0 = 0 dvtp1 = 0
+ dvt0 = 4.4955 dvt1 = 0.294 dvt2 = 0.015
+ dvt0w = -4.9772 dvt1w = 1.1472E6 dvt2w = -8.96E-3
+ vfbsdoff = 0 u0 = -8.087662470994137E-3 lu0 = 5.089322996095522E-8
+ wu0 = 6.400768948190965E-9 pu0 = -2.054378768474559E-14 ua = -1.780089536958452E-9
+ lua = 2.961634112431795E-15 wua = 3.822425751496523E-16 pua = -1.113971342228192E-21
+ ub = -9.594339868352658E-19 lub = 6.345627907651832E-24 wub = 6.679247348413641E-25
+ pub = -2.721782827104427E-30 uc = -5.744470591310368E-11 luc = 4.173698566665478E-17
+ wuc = -1.155804339358868E-17 puc = -8.650605684295114E-24 ud = 0
+ up = 0 lp = 1 eu = 1.67
+ vsat = 2.256235247288263E5 lvsat = -0.500138211986416 wvsat = -0.077971522843417
+ pvsat = 2.159823604784876E-7 a0 = 1.523261092041923 la0 = -1.352166277157789E-6
+ wa0 = -1.006178367357374E-7 pa0 = 5.355278105153723E-13 ags = -0.694088580084904
+ lags = 3.849340929179923E-6 wags = 3.141241013755496E-7 pags = -1.324634279476367E-12
+ b0 = 5.748989788328406E-7 lb0 = -1.785060546010789E-12 wb0 = -2.49020715441161E-13
+ pb0 = 7.554312541054479E-19 b1 = 1.748827207062223E-9 lb1 = -6.673801520849888E-15
+ wb1 = -8.952589012762618E-16 pb1 = 3.738440097574304E-21 keta = 0.054538012499851
+ lketa = -1.692828002930574E-7 wketa = -1.48471278339067E-8 pketa = 5.576678684112925E-14
+ a1 = 0 a2 = 0.8 rdsw = 547.88
+ rdswmin = 0 rdw = 0 rdwmin = 0
+ rsw = 0 rswmin = 0 prwb = -0.32348
+ prwg = 0.1376 wr = 1 voff = -5.726465037844519E-3
+ lvoff = -6.698474920590973E-7 wvoff = -1.013531957002558E-7 pvoff = 2.87672975737006E-13
+ voffl = 0 minv = 0 nfactor = 1.87556588426301
+ lnfactor = 7.612559286236414E-7 wnfactor = -9.937129857125158E-9 pnfactor = -2.51529652589471E-13
+ eta0 = 0.160612523 leta0 = -3.24706275293724E-7 etab = -0.140472583
+ letab = 2.83862718653004E-7 dsub = 0.8641982 ldsub = -1.2253066992216E-6
+ cit = 2.559200769230768E-5 wcit = -8.347839300801534E-12 cdsc = 1.3E-4
+ cdscb = 7.8E-4 cdscd = 0 pclm = 0.096180572127583
+ lpclm = -1.453741581280999E-6 wpclm = 2.164043750898719E-7 ppclm = 5.614831803240171E-13
+ pdiblc1 = 0.39 pdiblc2 = 3.257234435174975E-3 lpdiblc2 = -1.225021668976709E-8
+ wpdiblc2 = -1.437077639938094E-9 ppdiblc2 = 6.25012004084831E-15 pdiblcb = -1.060206889918154
+ lpdiblcb = 3.364203330107643E-6 wpdiblcb = 3.385863585590781E-7 ppdiblcb = -1.363821789239664E-12
+ drout = 0.56 pscbe1 = 8.782554376506895E8 lpscbe1 = -158.7010884903466
+ wpscbe1 = -41.89735092576551 ppscbe1 = 8.496732490924136E-5 pscbe2 = 9.97523101600994E-9
+ lpscbe2 = -4.214269800021436E-16 wpscbe2 = -1.841980030323081E-16 ppscbe2 = 1.138082006684697E-22
+ pvag = 0 delta = 0.01 fprout = 0
+ pdits = 0 pditsl = 0 pditsd = 0
+ lambda = 0 vtl = 0 lc = 5E-9
+ xn = 3 alpha0 = -4.670336219471758E-10 lalpha0 = 9.781661468692165E-16
+ walpha0 = 2.709775333198139E-16 palpha0 = -5.621175190688957E-22 alpha1 = -6.280417975398602E-10
+ lalpha1 = 1.273656984154662E-15 walpha1 = 3.362489918413185E-16 palpha1 = -6.819071996758843E-22
+ beta0 = 248.32066466536867 lbeta0 = -6.682575483712932E-4 wbeta0 = -1.090592651870975E-4
+ pbeta0 = 3.125891978992027E-10 aigbacc = 0.43 bigbacc = 0.054
+ cigbacc = 0.075 nigbacc = 1 aigbinv = 0.35
+ bigbinv = 0.03 cigbinv = 6E-3 eigbinv = 1.1
+ nigbinv = 3 aigc = 0.43 bigc = 0.054
+ cigc = 0.075 aigsd = 0.43 bigsd = 0.054
+ cigsd = 0.075 dlcig = 0 nigc = 1
+ poxedge = 1 pigcd = 1 ntox = 1
+ toxref = 4.23E-9 agidl = -3.70207214470676E-9 lagidl = 5.964385348251651E-15
+ wagidl = 1.898816556736782E-15 pagidl = -2.642324251166283E-21 bgidl = 3.667755206265639E9
+ lbgidl = -5.410175545244242E3 wbgidl = -1.081487152129481E3 pbgidl = 2.193242966672763E-3
+ cgidl = 300 egidl = 0.1 noia = 1.5E42
+ noib = 0 noic = 0 em = 4.1E7
+ af = 1 ef = 1 kf = 0
+ lintnoi = -2E-7 tnoia = 2.5E7 tnoib = 0
+ ntnoi = 1 rnoia = 0.69 rnoib = 0.34
+ xpart = 0 cgso = {5.248925E-11/sw_func_tox_lv_ratio} cgdo = {5.248925E-11/sw_func_tox_lv_ratio}
+ cgbo = {0/sw_func_tox_lv_ratio} ckappas = 0.6 cf = 1.2E-11
+ clc = 1E-7 cle = 0.6 dlc = -3E-9
+ dwc = 0 vfbcv = -0.14469 noff = 3.9
+ voffcv = -0.10701 acde = 0.8 moin = 18.13
+ cgsl = {9.548271750000001E-12/sw_func_tox_lv_ratio} cgdl = {9.548271750000001E-12/sw_func_tox_lv_ratio} ijthsrev = 0.1
+ ijthsfwd = 0.1 xjbvs = 1 bvs = 12.69
+ jss = 2.1483E-5 jsws = 8.040000000000001E-10 cjs = {sw_psd_nw_cj}
+ mjs = 0.34629 mjsws = 0.29781 cjsws = {9.888891999999999E-11*sw_func_psd_nw_cj}
+ cjswgs = {2.39155046E-10*sw_func_psd_nw_cj} mjswgs = 0.9274 pbs = 0.6587
+ pbsws = 0.7418 pbswgs = 1.4338 xrcrg1 = 12
+ xrcrg2 = 1 rbpb = 50 rbpd = 50
+ rbps = 50 rbdb = 50 rbsb = 50
+ gbmin = 1E-12 tnom = 30 ute = 2.529363131912557
+ lute = -8.045965072329673E-6 wute = -1.222418621672537E-6 pute = 2.992265988436588E-12
+ kt1 = -0.102613801415074 lkt1 = -1.008173900551745E-6 wkt1 = -1.023524896802801E-7
+ pkt1 = 3.259175391152226E-13 kt1l = 0 kt2 = -0.072913465892266
+ lkt2 = 1.727849784038291E-8 wkt2 = 7.144395745472675E-9 pkt2 = -7.004568252208077E-15
+ ua1 = 3.2341880759269E-9 lua1 = -6.452245610925686E-15 wua1 = -1.322701337288858E-15
+ pua1 = 2.615690043153508E-21 ub1 = -8.895285351350563E-19 lub1 = 1.562866224946815E-24
+ wub1 = 6.524514488709637E-25 pub1 = -6.335737772368842E-31 uc1 = -6.975765309212327E-10
+ luc1 = 1.522854089461196E-15 wuc1 = 3.005572528759538E-16 puc1 = -6.173531696056709E-22
+ at = 1.880571842102656E5 lat = -0.516915222869843 wat = -0.054646692967554
+ pat = 2.267469854036295E-7 prt = 0 njs = 1.3632
+ xtis = 5.2 tpb = 2.0386E-3 tpbsw = 1.246E-3
+ tpbswg = 0 tcj = 1.2407E-3 tcjsw = 3.7357E-4
+ tcjswg = 2E-12 tvoff = 0 tvfbsdoff = 0
+ saref = 3E-6 sbref = 3E-6 wlod = 0
+ ku0 = 4.5E-8 kvsat = 0.5 kvth0 = 3.29E-8
+ tku0 = 0 llodku0 = 0 wlodku0 = 1
+ llodvth = 0 wlodvth = 1 lku0 = 0
+ wku0 = 2.5E-7 pku0 = 0 lkvth0 = 0
+ wkvth0 = 2E-7 pkvth0 = 0 stk2 = 0
+ lodk2 = 1 steta0 = 0 lodeta0 = 1

.model pshort_model.44 pmos
+ level = 54 lmin = 1E-6 lmax = 2E-6 wmin = 4.2E-7
+ wmax = 5.5E-7 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 4.23E-9
+ toxm = 4.23E-9 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 9.999999999999999E22 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {7.3039E-9+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {-1.3994E-8-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = -5.722E-9 dwb = -1.7864E-8 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = -1.239560168718978 lvth0 = 3.49584260157244E-7
+ wvth0 = 8.765882778689792E-8 pvth0 = -1.530419221276315E-13 k1 = 0.307608382905938
+ lk1 = 3.097804817031309E-7 wk1 = 5.637497184102616E-8 pk1 = -1.26193965491908E-13
+ k2 = -0.01356698733887 lk2 = -2.131421374876534E-8 wk2 = 1.610867521918389E-8
+ pk2 = 2.856707318427954E-15 k3 = -15.845 k3b = 2
+ w0 = 0 lpe0 = 0 lpeb = 0
+ vbm = -3 dvtp0 = 0 dvtp1 = 0
+ dvt0 = 4.4955 dvt1 = 0.294 dvt2 = 0.015
+ dvt0w = -4.9772 dvt1w = 1.1472E6 dvt2w = -8.96E-3
+ vfbsdoff = 0 u0 = 0.036230221465893 lu0 = -3.898290684844382E-8
+ wu0 = -1.150063072032428E-8 pu0 = 1.576003602620731E-14 ua = 2.567292475339789E-9
+ lua = -5.854804439924891E-15 wua = -1.139336278387099E-15 pua = 1.971772313798097E-21
+ ub = 1.9374185703351E-18 lub = 4.708456839410171E-25 wub = -8.857999929658755E-25
+ pub = 4.291522761919218E-31 uc = -1.113855137859757E-10 luc = 1.511282967431447E-16
+ wuc = 1.302836111896586E-18 puc = -3.473231499086517E-23 ud = 0
+ up = 0 lp = 1 eu = 1.67
+ vsat = -2.519341898637795E5 lvsat = 0.468343102514813 wvsat = 0.122274876534341
+ pvsat = -1.90114934502814E-7 a0 = -0.460648598564659 la0 = 2.671178768476072E-6
+ wa0 = 8.358438698615909E-7 pa0 = -1.36360529292353E-12 ags = 2.566346127041278
+ lags = -2.762781531655489E-6 wags = -1.002939871576192E-6 pags = 1.34635565290209E-12
+ b0 = -5.806454793196655E-7 lb0 = 5.583697485889957E-13 wb0 = 2.513058400336807E-13
+ pb0 = -2.592249964788655E-19 b1 = 1.814970867759266E-10 lb1 = -3.495274844870722E-15
+ wb1 = 1.79030382252129E-16 pb1 = 1.559794322050129E-21 keta = -0.086578017721592
+ lketa = 1.168988156036661E-7 wketa = 4.02663601774111E-8 pketa = -5.600270548396712E-14
+ a1 = 0 a2 = 2.493466944287999 la2 = -3.434330641412732E-6
+ wa2 = -6.865182901721894E-7 pa2 = 1.392250854249718E-12 rdsw = 547.88
+ rdswmin = 0 rdw = 0 rdwmin = 0
+ rsw = 0 rswmin = 0 prwb = -0.32348
+ prwg = 0.1376 wr = 1 voff = -0.505117774979488
+ lvoff = 3.429120918068368E-7 wvoff = 1.347027094235455E-7 pvoff = -1.910455671832015E-13
+ voffl = 0 minv = 0 nfactor = 3.162330256221784
+ lnfactor = -1.84828677653629E-6 wnfactor = -3.935630573398819E-7 pnfactor = 5.264591248344299E-13
+ eta0 = -0.502700126 leta0 = 1.020483817126488E-6 etab = -0.0958645212594
+ letab = 1.933981047398076E-7 wetab = 1.41594397348014E-7 petab = -2.871517386890042E-13
+ dsub = 0.26 cit = 2.559200769230768E-5 wcit = -8.347839300801534E-12
+ cdsc = 1.3E-4 cdscb = 7.8E-4 cdscd = 0
+ pclm = -2.104065365293126 lpclm = 3.00833077685695E-6 wpclm = 1.079745749308069E-6
+ ppclm = -1.189362766493997E-12 pdiblc1 = 0.377007194731406 lpdiblc1 = 2.63492531710462E-8
+ wpdiblc1 = 6.676407534881793E-9 ppdiblc1 = -1.353967436384986E-14 pdiblc2 = -6.086619182045466E-3
+ lpdiblc2 = 6.699006319712552E-9 wpdiblc2 = 3.335743831985534E-9 ppdiblc2 = -3.429104630355145E-15
+ pdiblcb = 1.445413779836307 lpdiblcb = -1.717165320706365E-6 wpdiblcb = -6.77172717118156E-7
+ ppdiblcb = 6.961254271248588E-13 drout = -0.248320924845186 ldrout = 1.639265135734939E-6
+ wdrout = 2.520414255450013E-7 pdrout = -5.111369865081561E-13 pscbe1 = 7.294316563678579E8
+ lpscbe1 = 143.11175406586042 wpscbe1 = 38.444234753608896 ppscbe1 = -7.79644467495018E-5
+ pscbe2 = 1.067411972222421E-8 lpscbe2 = -1.838764889540216E-15 wpscbe2 = -3.26965637042095E-16
+ ppscbe2 = 4.033392492287095E-22 pvag = 0 delta = 0.01
+ fprout = 0 pdits = 0 pditsl = 0
+ pditsd = 0 lambda = 0 vtl = 0
+ lc = 5E-9 xn = 3 alpha0 = -7.177123403619283E-11
+ lalpha0 = 1.765787673343978E-16 walpha0 = -1.25783332267129E-17 palpha0 = 1.293037561706214E-23
+ alpha1 = -1.028030447546043E-10 lalpha1 = 2.084790963711962E-16 walpha1 = 1.720790407508544E-21
+ palpha1 = -1.768951889433893E-27 beta0 = -177.84630437561194 lbeta0 = 1.96003950840187E-4
+ wbeta0 = 9.411334218787833E-5 pbeta0 = -9.944241178595994E-11 aigbacc = 0.43
+ bigbacc = 0.054 cigbacc = 0.075 nigbacc = 1
+ aigbinv = 0.35 bigbinv = 0.03 cigbinv = 6E-3
+ eigbinv = 1.1 nigbinv = 3 aigc = 0.43
+ bigc = 0.054 cigc = 0.075 aigsd = 0.43
+ bigsd = 0.054 cigsd = 0.075 dlcig = 0
+ nigc = 1 poxedge = 1 pigcd = 1
+ ntox = 1 toxref = 4.23E-9 agidl = 4.777018223142507E-10
+ lagidl = -2.512146099579354E-15 wagidl = -2.203457107813246E-16 pagidl = 1.655311397413228E-21
+ bgidl = 1E9 cgidl = 300 egidl = 0.1
+ noia = 1.5E42 noib = 0 noic = 0
+ em = 4.1E7 af = 1 ef = 1
+ kf = 0 lintnoi = -2E-7 tnoia = 2.5E7
+ tnoib = 0 ntnoi = 1 rnoia = 0.69
+ rnoib = 0.34 xpart = 0 cgso = {5.248925E-11/sw_func_tox_lv_ratio}
+ cgdo = {5.248925E-11/sw_func_tox_lv_ratio} cgbo = {0/sw_func_tox_lv_ratio} ckappas = 0.6
+ cf = 1.2E-11 clc = 1E-7 cle = 0.6
+ dlc = -3E-9 dwc = 0 vfbcv = -0.14469
+ noff = 3.9 voffcv = -0.10701 acde = 0.8
+ moin = 18.13 cgsl = {9.548271750000001E-12/sw_func_tox_lv_ratio} cgdl = {9.548271750000001E-12/sw_func_tox_lv_ratio}
+ ijthsrev = 0.1 ijthsfwd = 0.1 xjbvs = 1
+ bvs = 12.69 jss = 2.1483E-5 jsws = 8.040000000000001E-10
+ cjs = {sw_psd_nw_cj} mjs = 0.34629 mjsws = 0.29781
+ cjsws = {9.888891999999999E-11*sw_func_psd_nw_cj} cjswgs = {2.39155046E-10*sw_func_psd_nw_cj} mjswgs = 0.9274
+ pbs = 0.6587 pbsws = 0.7418 pbswgs = 1.4338
+ xrcrg1 = 12 xrcrg2 = 1 rbpb = 50
+ rbpd = 50 rbps = 50 rbdb = 50
+ rbsb = 50 gbmin = 1E-12 tnom = 30
+ ute = -4.487892038661162 lute = 6.184944206531783E-6 wute = 1.453818917647113E-6
+ pute = -2.435111626453191E-12 kt1 = -0.592176172339095 lkt1 = -1.534728706628089E-8
+ wkt1 = 6.966019560109429E-8 pkt1 = -2.292212248318126E-14 kt1l = 0
+ kt2 = -0.079096994455688 lkt2 = 2.981861956466084E-8 wkt2 = 1.278420991362158E-8
+ pkt2 = -1.844204370744404E-14 ua1 = -4.54665601797395E-9 lua1 = 9.32721284137611E-15
+ wua1 = 1.872467236318508E-15 pua1 = -3.864073482099346E-21 ub1 = 4.457726949489547E-18
+ lub1 = -9.281303730806067E-24 wub1 = -1.55832219889895E-24 pub1 = 3.849848651156727E-30
+ uc1 = 2.078721194950896E-10 luc1 = -3.133849081993009E-16 wuc1 = -5.977362524585615E-17
+ puc1 = 1.133935272548221E-22 at = -2.518398514602474E5 lat = 0.375190686705529
+ wat = 0.13812256570444 pat = -1.641867579520692E-7 prt = 0
+ njs = 1.3632 xtis = 5.2 tpb = 2.0386E-3
+ tpbsw = 1.246E-3 tpbswg = 0 tcj = 1.2407E-3
+ tcjsw = 3.7357E-4 tcjswg = 2E-12 tvoff = 0
+ tvfbsdoff = 0 saref = 3E-6 sbref = 3E-6
+ wlod = 0 ku0 = 4.5E-8 kvsat = 0.5
+ kvth0 = 3.29E-8 tku0 = 0 llodku0 = 0
+ wlodku0 = 1 llodvth = 0 wlodvth = 1
+ lku0 = 0 wku0 = 2.5E-7 pku0 = 0
+ lkvth0 = 0 wkvth0 = 2E-7 pkvth0 = 0
+ stk2 = 0 lodk2 = 1 steta0 = 0
+ lodeta0 = 1

.model pshort_model.45 pmos
+ level = 54 lmin = 5E-7 lmax = 1E-6 wmin = 4.2E-7
+ wmax = 5.5E-7 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 4.23E-9
+ toxm = 4.23E-9 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 9.999999999999999E22 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {7.3039E-9+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {-1.3994E-8-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = -5.722E-9 dwb = -1.7864E-8 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = -0.889557183849071 lvth0 = -1.021460825320138E-8
+ wvth0 = -7.91290474468747E-8 pvth0 = 1.841401215818394E-14 k1 = 0.603238458959026
+ lk1 = 5.876311081469773E-9 wk1 = -9.255817820667973E-8 pk1 = 2.690752555933306E-14
+ k2 = -0.028876062754494 lk2 = -5.576667930409036E-9 wk2 = 2.466582728351857E-8
+ pk2 = -5.939942317883322E-15 k3 = -15.845 k3b = 2
+ w0 = 0 lpe0 = 0 lpeb = 0
+ vbm = -3 dvtp0 = 0 dvtp1 = 0
+ dvt0 = 4.4955 dvt1 = 0.294 dvt2 = 0.015
+ dvt0w = -4.9772 dvt1w = 1.1472E6 dvt2w = -8.96E-3
+ vfbsdoff = 0 u0 = -6.026822870679344E-3 lu0 = 4.456827645020098E-9
+ wu0 = 6.434132125885552E-9 pu0 = -2.676684962542244E-15 ua = -3.974434941427992E-9
+ lua = 8.700128437833872E-16 wua = 1.307726813275027E-15 pua = -5.437791796734684E-22
+ ub = 2.771191594984537E-18 lub = -3.862629801223088E-25 wub = -7.538101162414936E-25
+ pub = 2.934682667977778E-31 uc = 5.71460387077808E-11 luc = -2.212011684180702E-17
+ wuc = -5.076442109647627E-17 puc = 1.879220061225562E-23 ud = 0
+ up = 0 lp = 1 eu = 1.67
+ vsat = 2.853199072152592E5 lvsat = -0.083947662233274 wvsat = -0.108264698191764
+ pvsat = 4.687698184072578E-8 a0 = 3.631506692597601 la0 = -1.535507764975236E-6
+ wa0 = -1.224091978408693E-6 pa0 = 7.539840398681428E-13 ags = 0.209281556720716
+ lags = -3.397474381407945E-7 wags = -8.601798644322097E-8 pags = 4.037709580480172E-13
+ b0 = 7.611794495848625E-8 lb0 = -1.167751704078529E-13 wb0 = -4.52085924163266E-14
+ pb0 = 4.558828190655263E-20 b1 = 6.625365667570082E-9 lb1 = -1.011949441950415E-14
+ wb1 = -3.789755594648544E-15 pb1 = 5.639658680872299E-21 keta = -0.012990877802709
+ lketa = 4.125211881273271E-8 wketa = 1.280859263004662E-8 pketa = -2.777644993848701E-14
+ a1 = 0 a2 = -2.586933888575998 la2 = 1.788260449961464E-6
+ wa2 = 1.373036580344379E-6 pa2 = -7.249468379828676E-13 rdsw = 547.88
+ rdswmin = 0 rdw = 0 rdwmin = 0
+ rsw = 0 rswmin = 0 prwb = -0.32348
+ prwg = 0.1376 wr = 1 voff = -0.17839027328982
+ lvoff = 7.04014079987785E-9 wvoff = -5.540932600455387E-8 pvoff = 4.387323892459496E-15
+ voffl = 0 minv = 0 nfactor = 0.856087110130422
+ lnfactor = 5.225035027278776E-7 wnfactor = 1.751534573522464E-7 pnfactor = -5.817462767090155E-14
+ eta0 = 0.49 etab = 0.189717944859996 letab = -1.001772434413381E-7
+ wetab = -2.83194304144749E-7 petab = 1.495259489811382E-13 dsub = 0.349430903910948
+ ldsub = -9.193389604960754E-8 wdsub = -6.91651784867768E-8 pdsub = 7.110097350226472E-14
+ cit = 4.205679360719998E-5 lcit = -1.69256023430783E-11 wcit = -1.716295725430473E-11
+ pcit = 9.061835474785846E-18 cdsc = 1.3E-4 cdscb = 7.8E-4
+ cdscd = 0 pclm = 1.107998999936059 lpclm = -2.936328458262686E-7
+ wpclm = -2.033710565736464E-7 ppclm = 1.296659125507364E-13 pdiblc1 = 1.130784855108158
+ lpdiblc1 = -7.48525136364331E-7 wpdiblc1 = -2.864685469621054E-7 ppdiblc1 = 2.87809821119599E-13
+ pdiblc2 = 2.84137468502792E-3 lpdiblc2 = -2.478864239712482E-9 wpdiblc2 = -1.577370612891632E-9
+ ppdiblc2 = 1.621518061605244E-15 pdiblcb = 0.433591436595692 lpdiblcb = -6.770240937231319E-7
+ wpdiblcb = -3.526047181401279E-7 ppdiblcb = 3.624734189914338E-13 drout = 1.961888928147833
+ ldrout = -6.328040706236494E-7 wdrout = -5.447987702123717E-7 pdrout = 3.080051726480743E-13
+ pscbe1 = 9.411366872642841E8 lpscbe1 = -74.51847723529477 wpscbe1 = -76.8884695072178
+ ppscbe1 = 4.059618923817691E-5 pscbe2 = 4.451265140061979E-8 lpscbe2 = -3.662436939255074E-14
+ wpscbe2 = -1.448198864728779E-14 ppscbe2 = 1.495453304348517E-20 pvag = 0
+ delta = 0.01 fprout = 0 pdits = 0
+ pditsl = 0 pditsd = 0 lambda = 0
+ vtl = 0 lc = 5E-9 xn = 3
+ alpha0 = 1E-10 alpha1 = 1E-10 beta0 = 17.597724801275803
+ lbeta0 = -4.910165825303411E-6 wbeta0 = -5.820293565556012E-6 pbeta0 = 3.288166564941516E-12
+ aigbacc = 0.43 bigbacc = 0.054 cigbacc = 0.075
+ nigbacc = 1 aigbinv = 0.35 bigbinv = 0.03
+ cigbinv = 6E-3 eigbinv = 1.1 nigbinv = 3
+ aigc = 0.43 bigc = 0.054 cigc = 0.075
+ aigsd = 0.43 bigsd = 0.054 cigsd = 0.075
+ dlcig = 0 nigc = 1 poxedge = 1
+ pigcd = 1 ntox = 1 toxref = 4.23E-9
+ agidl = -3.286037564875388E-9 lagidl = 1.356932825578949E-15 wagidl = 2.267089122473683E-15
+ pagidl = -9.017417619549217E-22 bgidl = 1E9 cgidl = 300
+ egidl = 0.1 noia = 1.5E42 noib = 0
+ noic = 0 em = 4.1E7 af = 1
+ ef = 1 kf = 0 lintnoi = -2E-7
+ tnoia = 2.5E7 tnoib = 0 ntnoi = 1
+ rnoia = 0.69 rnoib = 0.34 xpart = 0
+ cgso = {5.248925E-11/sw_func_tox_lv_ratio} cgdo = {5.248925E-11/sw_func_tox_lv_ratio} cgbo = {0/sw_func_tox_lv_ratio}
+ ckappas = 0.6 cf = 1.2E-11 clc = 1E-7
+ cle = 0.6 dlc = -3E-9 dwc = 0
+ vfbcv = -0.14469 noff = 3.9 voffcv = -0.10701
+ acde = 0.8 moin = 18.13 cgsl = {9.548271750000001E-12/sw_func_tox_lv_ratio}
+ cgdl = {9.548271750000001E-12/sw_func_tox_lv_ratio} ijthsrev = 0.1 ijthsfwd = 0.1
+ xjbvs = 1 bvs = 12.69 jss = 2.1483E-5
+ jsws = 8.040000000000001E-10 cjs = {sw_psd_nw_cj} mjs = 0.34629
+ mjsws = 0.29781 cjsws = {9.888891999999999E-11*sw_func_psd_nw_cj} cjswgs = {2.39155046E-10*sw_func_psd_nw_cj}
+ mjswgs = 0.9274 pbs = 0.6587 pbsws = 0.7418
+ pbswgs = 1.4338 xrcrg1 = 12 xrcrg2 = 1
+ rbpb = 50 rbpd = 50 rbps = 50
+ rbdb = 50 rbsb = 50 gbmin = 1E-12
+ tnom = 30 ute = 3.070934721587373 lute = -1.585438997082587E-6
+ wute = -1.790657558259555E-6 pute = 9.001712570611535E-13 kt1 = -0.710280397833605
+ lkt1 = 1.060624394913696E-7 wkt1 = 9.737544534479292E-8 pkt1 = -5.141306663670652E-14
+ kt1l = 0 kt2 = -0.095347290823325 lkt2 = 4.652372922703586E-8
+ wkt2 = 2.805247054900079E-8 pkt2 = -3.413763242148625E-14 ua1 = 9.244178359835554E-9
+ lua1 = -4.849599408999524E-15 wua1 = -4.021609671814125E-15 pua1 = 2.194966850538102E-21
+ ub1 = -9.949121009685252E-18 lub1 = 5.52876308905012E-24 wub1 = 4.52142336364696E-24
+ pub1 = -2.400056830193718E-30 uc1 = -2.250710639675656E-10 luc1 = 1.31675489082107E-16
+ wuc1 = 1.038939155711698E-16 puc1 = -5.485474069459082E-23 at = 1.200789958563693E5
+ lat = -7.137425309784661E-3 wat = -0.021408771158242 pat = -1.904580332748519E-10
+ prt = 0 njs = 1.3632 xtis = 5.2
+ tpb = 2.0386E-3 tpbsw = 1.246E-3 tpbswg = 0
+ tcj = 1.2407E-3 tcjsw = 3.7357E-4 tcjswg = 2E-12
+ tvoff = 0 tvfbsdoff = 0 saref = 2.75E-6
+ sbref = 2.74E-6 wlod = 0 ku0 = 4.5E-8
+ kvsat = 0.5 kvth0 = 3.29E-8 tku0 = 0
+ llodku0 = 0 wlodku0 = 1 llodvth = 0
+ wlodvth = 1 lku0 = 0 wku0 = 2.5E-7
+ pku0 = 0 lkvth0 = 0 wkvth0 = 2E-7
+ pkvth0 = 0 stk2 = 0 lodk2 = 1
+ steta0 = 0 lodeta0 = 1

.model pshort_model.46 pmos
+ level = 54 lmin = 2.5E-7 lmax = 5E-7 wmin = 4.2E-7
+ wmax = 5.5E-7 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 4.23E-9
+ toxm = 4.23E-9 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 9.999999999999999E22 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {7.3039E-9+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {-1.3994E-8-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = -5.722E-9 dwb = -1.7864E-8 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = -0.724921142726069 lvth0 = -9.714046233365291E-8
+ wvth0 = -1.277573003613919E-7 pvth0 = 4.408914615801404E-14 k1 = -0.900993997288542
+ lk1 = 8.000929971907101E-7 wk1 = 3.605878914026057E-7 pk1 = -2.123481614415343E-13
+ k2 = 0.526751257650574 lk2 = -2.989412255764399E-7 wk2 = -1.308646732158936E-7
+ pk2 = 7.617829557980033E-14 k3 = -15.845 k3b = 2
+ w0 = 0 lpe0 = 0 lpeb = 0
+ vbm = -3 dvtp0 = 0 dvtp1 = 0
+ dvt0 = 4.4955 dvt1 = 0.294 dvt2 = 0.015
+ dvt0w = -4.9772 dvt1w = 1.1472E6 dvt2w = -8.96E-3
+ vfbsdoff = 0 u0 = 3.020883555092865E-3 lu0 = -3.202527753105184E-10
+ wu0 = 2.440701745045986E-9 pu0 = -5.682016426235236E-16 ua = -1.845128543170706E-9
+ lua = -2.5423538281968E-16 wua = 4.51209123688069E-16 pua = -9.15481177838299E-23
+ ub = 1.262665005043841E-18 lub = 4.102209570472993E-25 wub = -2.16749066432308E-25
+ pub = 9.906477231125612E-33 uc = 3.174719976618334E-11 luc = -8.709834666710863E-18
+ wuc = -3.188988615903592E-17 puc = 8.82667265970637E-24 ud = 0
+ up = 0 lp = 1 eu = 1.67
+ vsat = 2.505617809829932E5 lvsat = -0.065595788680152 wvsat = -0.088203669306049
+ pvsat = 3.628499932141457E-8 a0 = 3.081493447238975 la0 = -1.245107371584827E-6
+ wa0 = -7.855744731388738E-7 pa0 = 5.224520592957413E-13 ags = -5.169102667468366
+ lags = 2.499974891620349E-6 wags = 2.593717549462944E-6 pags = -1.011097248084007E-12
+ b0 = -6.93228503957029E-7 lb0 = 2.894305224621521E-13 wb0 = 2.77967736428662E-13
+ pb0 = -1.250449416076551E-19 b1 = -1.297555208189485E-8 lb1 = 2.295549412003433E-16
+ wb1 = 5.820117609421236E-15 pb1 = 5.65760947601904E-22 keta = 0.461380709274354
+ lketa = -2.092103867049112E-7 wketa = -2.425398300426632E-7 pketa = 1.070444530516317E-13
+ a1 = 0 a2 = 0.344390971874074 la2 = 2.405560995421513E-7
+ wa2 = 2.439295199082013E-7 pa2 = -1.287918593572914E-13 rdsw = 547.88
+ rdswmin = 0 rdw = 0 rdwmin = 0
+ rsw = 0 rswmin = 0 prwb = -0.32348
+ prwg = 0.1376 wr = 1 voff = 0.121110876437984
+ lvoff = -1.510928722426056E-7 wvoff = -1.222016589763966E-7 pvoff = 3.965287419359678E-14
+ voffl = 0 minv = 0 nfactor = -0.858849054115481
+ lnfactor = 1.427969218215743E-6 wnfactor = 9.560064352837215E-7 pnfactor = -4.704556297829852E-13
+ eta0 = 0.641016265880455 leta0 = -7.973477618968965E-8 weta0 = 1.039134039451698E-7
+ peta0 = -5.486503032220232E-14 etab = -0.240779022673171 letab = 1.271199894525635E-7
+ wetab = 1.421838050314795E-7 petab = -7.506858812660033E-14 dsub = 0.084956409252972
+ ldsub = 4.77054634358677E-8 wdsub = 1.362861133337624E-7 pdsub = -3.737484316347813E-14
+ cit = 1E-5 cdsc = 1.3E-4 cdscb = 7.8E-4
+ cdscd = 0 pclm = 0.508227799302933 lpclm = 2.303915085361421E-8
+ wpclm = 7.343079016828642E-8 ppclm = -1.648214090684319E-14 pdiblc1 = -0.834041556376561
+ lpdiblc1 = 2.888796309826629E-7 wpdiblc1 = 5.624527674555115E-7 ppdiblc1 = -1.604104458371296E-13
+ pdiblc2 = -8.832399647592394E-3 lpdiblc2 = 3.684748522619052E-9 wpdiblc2 = 3.623969715889701E-9
+ ppdiblc2 = -1.124727215907355E-15 pdiblcb = -1.448932269270644 lpdiblcb = 3.169258326898229E-7
+ wpdiblcb = 5.659842261596425E-7 ppdiblcb = -1.225305205315133E-13 drout = 0.500246963085075
+ ldrout = 1.389253472259061E-7 wdrout = 8.143183824473838E-8 pdrout = -2.263707384997834E-14
+ pscbe1 = 8E8 pscbe2 = -9.207670391416775E-8 lpscbe2 = 3.549317114139331E-14
+ wpscbe2 = 4.483067980303004E-14 ppscbe2 = -1.636184414626125E-20 pvag = 0
+ delta = 0.01 fprout = 0 pdits = 0
+ pditsl = 0 pditsd = 0 lambda = 0
+ vtl = 0 lc = 5E-9 xn = 3
+ alpha0 = 1E-10 alpha1 = 1E-10 beta0 = 11.031865078662536
+ lbeta0 = -1.443470682080276E-6 wbeta0 = -2.830961704369924E-7 pbeta0 = 3.645927866874142E-13
+ aigbacc = 0.43 bigbacc = 0.054 cigbacc = 0.075
+ nigbacc = 1 aigbinv = 0.35 bigbinv = 0.03
+ cigbinv = 6E-3 eigbinv = 1.1 nigbinv = 3
+ aigc = 0.43 bigc = 0.054 cigc = 0.075
+ aigsd = 0.43 bigsd = 0.054 cigsd = 0.075
+ dlcig = 0 nigc = 1 poxedge = 1
+ pigcd = 1 ntox = 1 toxref = 4.23E-9
+ agidl = 7.56094694422565E-9 lagidl = -4.37014483141229E-15 wagidl = -4.577744995040359E-15
+ pagidl = 2.712248514083082E-21 bgidl = 1E9 cgidl = 300
+ egidl = 0.1 noia = 1.5E42 noib = 0
+ noic = 0 em = 4.1E7 af = 1
+ ef = 1 kf = 0 lintnoi = -2E-7
+ tnoia = 2.5E7 tnoib = 0 ntnoi = 1
+ rnoia = 0.69 rnoib = 0.34 xpart = 0
+ cgso = {5.248925E-11/sw_func_tox_lv_ratio} cgdo = {5.248925E-11/sw_func_tox_lv_ratio} cgbo = {0/sw_func_tox_lv_ratio}
+ ckappas = 0.6 cf = 1.2E-11 clc = 1E-7
+ cle = 0.6 dlc = -3E-9 dwc = 0
+ vfbcv = -0.14469 noff = 3.9 voffcv = -0.10701
+ acde = 0.8 moin = 18.13 cgsl = {9.548271750000001E-12/sw_func_tox_lv_ratio}
+ cgdl = {9.548271750000001E-12/sw_func_tox_lv_ratio} ijthsrev = 0.1 ijthsfwd = 0.1
+ xjbvs = 1 bvs = 12.69 jss = 2.1483E-5
+ jsws = 8.040000000000001E-10 cjs = {sw_psd_nw_cj} mjs = 0.34629
+ mjsws = 0.29781 cjsws = {9.888891999999999E-11*sw_func_psd_nw_cj} cjswgs = {2.39155046E-10*sw_func_psd_nw_cj}
+ mjswgs = 0.9274 pbs = 0.6587 pbsws = 0.7418
+ pbswgs = 1.4338 xrcrg1 = 12 xrcrg2 = 1
+ rbpb = 50 rbpd = 50 rbps = 50
+ rbdb = 50 rbsb = 50 gbmin = 1E-12
+ tnom = 30 ute = -0.314182380844868 lute = 2.018622115964068E-7
+ wute = 6.416169989237528E-8 pute = -7.915105341196787E-14 kt1 = -0.292991013960416
+ lkt1 = -1.142613477210677E-7 wkt1 = -3.670259618093396E-8 pkt1 = 1.937853035237896E-14
+ kt1l = 0 kt2 = 0.11816025535924 lkt2 = -6.620569306680429E-8
+ wkt2 = -7.730505840504167E-8 pkt2 = 2.148987857590073E-14 ua1 = 6.47145047960312E-12
+ lua1 = 2.77989866575051E-17 wua1 = 2.597988990786305E-16 pua1 = -6.556549799042145E-23
+ ub1 = 6.886285482736941E-19 lub1 = -8.784102455750771E-26 wub1 = -5.119820507394646E-26
+ pub1 = 1.423248663209623E-32 uc1 = 2.29278426924414E-11 luc1 = 7.350423525032491E-19
+ wuc1 = 5.643697136572567E-19 puc1 = -2.979804363744676E-25 at = 2.865015407589461E5
+ lat = -0.095006531947806 wat = -0.113795175282545 pat = 4.85884547075077E-8
+ prt = 0 njs = 1.3632 xtis = 5.2
+ tpb = 2.0386E-3 tpbsw = 1.246E-3 tpbswg = 0
+ tcj = 1.2407E-3 tcjsw = 3.7357E-4 tcjswg = 2E-12
+ tvoff = 0 tvfbsdoff = 0 saref = 1.75E-6
+ sbref = 1.74E-6 wlod = 0 ku0 = 4.5E-8
+ kvsat = 0.5 kvth0 = 3.29E-8 tku0 = 0
+ llodku0 = 0 wlodku0 = 1 llodvth = 0
+ wlodvth = 1 lku0 = 0 wku0 = 2.5E-7
+ pku0 = 0 lkvth0 = 0 wkvth0 = 2E-7
+ pkvth0 = 0 stk2 = 0 lodk2 = 1
+ steta0 = 0 lodeta0 = 1

.model pshort_model.47 pmos
+ level = 54 lmin = 1.8E-7 lmax = 2.5E-7 wmin = 4.2E-7
+ wmax = 5.5E-7 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 4.23E-9
+ toxm = 4.23E-9 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 9.999999999999999E22 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {7.3039E-9+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {-1.3994E-8-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = -5.722E-9 dwb = -1.7864E-8 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = -1.074362350021538 wvth0 = 3.084359664860149E-8
+ k1 = 1.9771626036824 wk1 = -4.032873889747282E-7 k2 = -0.548623310951092
+ wk2 = 1.431698015808613E-7 k3 = -15.845 k3b = 2
+ w0 = 0 lpe0 = 0 lpeb = 0
+ vbm = -3 dvtp0 = 0 dvtp1 = 0
+ dvt0 = 4.4955 dvt1 = 0.294 dvt2 = 0.015
+ dvt0w = -4.9772 dvt1w = 1.1472E6 dvt2w = -8.96E-3
+ vfbsdoff = 0 u0 = 1.86884542643077E-3 wu0 = 3.967227149312921E-10
+ ua = -2.759683785913846E-9 wua = 1.218851320631432E-16 ub = 2.738343656810462E-18
+ wub = -1.811127179887579E-25 uc = 4.155067912676367E-13 wuc = -1.378944913870628E-19
+ ud = 0 up = 0 lp = 1
+ eu = 1.67 vsat = 1.459552100000005E4 wvsat = 0.042323545255064
+ a0 = -1.39750338566326 wa0 = 1.093830606561477E-6 ags = 3.82400096153846
+ wags = -1.043479912600192E-6 b0 = 3.479334255584613E-7 wb0 = -1.718536285498808E-13
+ b1 = -1.214977923846153E-8 wb1 = 7.855316782054243E-15 keta = -0.291207124390809
+ wketa = 1.425287810183599E-7 a1 = 0 a2 = 1.209738035568015
+ wa2 = -2.193705482864379E-7 rdsw = 547.88 rdswmin = 0
+ rdw = 0 rdwmin = 0 rsw = 0
+ rswmin = 0 prwb = -0.32348 prwg = 0.1376
+ wr = 1 voff = -0.422412125427585 wvoff = 2.044073635576444E-8
+ voffl = 0 minv = 0 nfactor = 4.277952599969384
+ wnfactor = -7.363530542733283E-7 eta0 = 0.354188143120877 weta0 = -9.345133957686107E-8
+ etab = 0.216506865395968 wetab = -1.278587440231572E-7 dsub = 0.256566203329938
+ wdsub = 1.838427953536921E-9 cit = 1E-5 cdsc = 1.3E-4
+ cdscb = 7.8E-4 cdscd = 0 pclm = 0.591106020138416
+ wpclm = 1.413995420830546E-8 pdiblc1 = 0.205138663570569 wpdiblc1 = -1.458813300468691E-8
+ pdiblc2 = 4.422663601968923E-3 wpdiblc2 = -4.21986281877666E-10 pdiblcb = -0.308862076709012
+ wpdiblcb = 1.25207931745807E-7 drout = 1 pscbe1 = 8E8
+ pscbe2 = 3.560208488748307E-8 wpscbe2 = -1.402741531712351E-14 pvag = 0
+ delta = 0.01 fprout = 0 pdits = 0
+ pditsl = 0 pditsd = 0 lambda = 0
+ vtl = 0 lc = 5E-9 xn = 3
+ alpha0 = 1E-10 alpha1 = 1E-10 beta0 = 5.839300356155539
+ wbeta0 = 1.028445287062663E-6 aigbacc = 0.43 bigbacc = 0.054
+ cigbacc = 0.075 nigbacc = 1 aigbinv = 0.35
+ bigbinv = 0.03 cigbinv = 6E-3 eigbinv = 1.1
+ nigbinv = 3 aigc = 0.43 bigc = 0.054
+ cigc = 0.075 aigsd = 0.43 bigsd = 0.054
+ cigsd = 0.075 dlcig = 0 nigc = 1
+ poxedge = 1 pigcd = 1 ntox = 1
+ toxref = 4.23E-9 agidl = -8.159677080596609E-9 wagidl = 5.178965776946497E-15
+ bgidl = 1E9 cgidl = 300 egidl = 0.1
+ noia = 1.5E42 noib = 0 noic = 0
+ em = 4.1E7 af = 1 ef = 1
+ kf = 0 lintnoi = -2E-7 tnoia = 2.5E7
+ tnoib = 0 ntnoi = 1 rnoia = 0.69
+ rnoib = 0.34 xpart = 0 cgso = {5.248925E-11/sw_func_tox_lv_ratio}
+ cgdo = {5.248925E-11/sw_func_tox_lv_ratio} cgbo = {0/sw_func_tox_lv_ratio} ckappas = 0.6
+ cf = 1.2E-11 clc = 1E-7 cle = 0.6
+ dlc = -3E-9 dwc = 0 vfbcv = -0.14469
+ noff = 3.9 voffcv = -0.10701 acde = 0.8
+ moin = 18.13 cgsl = {9.548271750000001E-12/sw_func_tox_lv_ratio} cgdl = {9.548271750000001E-12/sw_func_tox_lv_ratio}
+ ijthsrev = 0.1 ijthsfwd = 0.1 xjbvs = 1
+ bvs = 12.69 jss = 2.1483E-5 jsws = 8.040000000000001E-10
+ cjs = {sw_psd_nw_cj} mjs = 0.34629 mjsws = 0.29781
+ cjsws = {9.888891999999999E-11*sw_func_psd_nw_cj} cjswgs = {2.39155046E-10*sw_func_psd_nw_cj} mjswgs = 0.9274
+ pbs = 0.6587 pbsws = 0.7418 pbswgs = 1.4338
+ xrcrg1 = 12 xrcrg2 = 1 rbpb = 50
+ rbpd = 50 rbps = 50 rbdb = 50
+ rbsb = 50 gbmin = 1E-12 tnom = 30
+ ute = 0.411972027246154 wute = -2.205666100057781E-7 kt1 = -0.704020798415384
+ wkt1 = 3.300735659536919E-8 kt1l = 0 kt2 = -0.12
+ ua1 = 1.064721219384616E-10 wua1 = 2.39416031146988E-17 ub1 = 3.7264E-19
+ uc1 = 2.557199406769231E-11 wuc1 = -5.075486294887338E-19 at = -5.526332660153837E4
+ wat = 0.060990983499516 prt = 0 njs = 1.3632
+ xtis = 5.2 tpb = 2.0386E-3 tpbsw = 1.246E-3
+ tpbswg = 0 tcj = 1.2407E-3 tcjsw = 3.7357E-4
+ tcjswg = 2E-12 tvoff = 0 tvfbsdoff = 0
+ saref = 1.1E-6 sbref = 1.1E-6 wlod = 0
+ ku0 = 4.5E-8 kvsat = 0.5 kvth0 = 3.29E-8
+ tku0 = 0 llodku0 = 0 wlodku0 = 1
+ llodvth = 0 wlodvth = 1 lku0 = 0
+ wku0 = 2.5E-7 pku0 = 0 lkvth0 = 0
+ wkvth0 = 2E-7 pkvth0 = 0 stk2 = 0
+ lodk2 = 1 steta0 = 0 lodeta0 = 1

.model pshort_model.48 pmos
+ level = 54 lmin = 1.5E-7 lmax = 1.8E-7 wmin = 4.2E-7
+ wmax = 5.5E-7 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 4.23E-9
+ toxm = 4.23E-9 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 9.999999999999999E22 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {7.3039E-9+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {-1.3994E-8-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = -5.722E-9 dwb = -1.7864E-8 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = -1.304407121733081 lvth0 = 4.784655197874038E-8
+ wvth0 = 1.540077730737422E-7 pvth0 = -2.561667072631217E-14 k1 = 2.817933506358009
+ lk1 = -1.748702585056946E-7 wk1 = -8.534295722542082E-7 pk1 = 9.362417241593253E-14
+ k2 = -1.151966695759153 lk2 = 1.254881839194589E-7 wk2 = 4.661951437286954E-7
+ pk2 = -6.718539486264373E-14 k3 = -15.845 k3b = 2
+ w0 = 0 lpe0 = 0 lpeb = 0
+ vbm = -3 dvtp0 = 0 dvtp1 = 0
+ dvt0 = 4.4955 dvt1 = 0.294 dvt2 = 0.015
+ dvt0w = -4.9772 dvt1w = 1.1472E6 dvt2w = -8.96E-3
+ vfbsdoff = 0 u0 = 1.77134374178224E-3 lu0 = 2.027918038667842E-11
+ wu0 = 4.489243563789747E-10 pu0 = -1.085731500142061E-17 ua = -3.214592974175342E-9
+ lua = 9.461565224813203E-17 wua = 3.654399631666797E-16 pua = -5.065648221156236E-23
+ ub = 4.237991721651763E-18 lub = -3.119088017102127E-25 wub = -9.840125946498852E-25
+ pub = 1.669935395469946E-31 uc = 3.196856017660247E-12 luc = -5.784872628989464E-19
+ wuc = -1.627007172673701E-18 puc = 3.097175683554453E-25 ud = 0
+ up = 0 lp = 1 eu = 1.67
+ vsat = 1.224579159717148E5 lvsat = -0.022434083805377 wvsat = -0.015425139686112
+ pvsat = 1.201103348354517E-8 a0 = -9.350451604330704 la0 = 1.654117794104204E-6
+ wa0 = 5.351777049839922E-6 pa0 = -8.856017648445972E-13 ags = 3.82400096153846
+ wags = -1.043479912600192E-6 b0 = 8.174586158830198E-7 lb0 = -9.765560528522431E-14
+ wb0 = -4.23233753153165E-13 pb0 = 5.228404935598788E-20 b1 = -9.699474615111789E-8
+ lb1 = 1.764673497822957E-14 wb1 = 5.328065027634854E-14 pb1 = -9.447924262811283E-21
+ keta = -1.180095644977254 lketa = 1.848781456197334E-7 wketa = 6.184327616098817E-7
+ pketa = -9.898231711526946E-14 a1 = 0 a2 = -1.125559225808243
+ la2 = 4.85713806799125E-7 wa2 = 1.030929390135772E-6 pa2 = -2.600473835925586E-13
+ rdsw = 547.88 rdswmin = 0 rdw = 0
+ rdwmin = 0 rsw = 0 rswmin = 0
+ prwb = -0.32348 prwg = 0.1376 wr = 1
+ voff = -0.59862190624913 lvoff = 3.664951989351158E-8 wvoff = 1.147820785713294E-7
+ pvoff = -1.962186708473093E-14 voffl = 0 minv = 0
+ nfactor = 14.389711705228454 lnfactor = -2.103124552784624E-6 wnfactor = -6.150110007508013E-6
+ pnfactor = 1.125996481189376E-12 eta0 = -0.50949905968053 leta0 = 1.79636573936259E-7
+ weta0 = 3.689600520428302E-7 peta0 = -9.617602052019636E-14 etab = 1.184185979311373
+ letab = -2.012656435450375E-7 wetab = -6.459465937163771E-7 petab = 1.077560556819934E-13
+ dsub = 0.236193716606241 ldsub = 4.237232768688309E-9 wdsub = 1.274569844000789E-8
+ pdsub = -2.268581373940125E-15 cit = 1E-5 cdsc = 1.3E-4
+ cdscb = 7.8E-4 cdscd = 0 pclm = 3.579253840500591
+ lpclm = -6.214988888614882E-7 wpclm = -1.585691081260605E-6 ppclm = 3.327456574051077E-13
+ pdiblc1 = 2.959952926744328 lpdiblc1 = -5.729683089689836E-7 wpdiblc1 = -1.489494201956665E-6
+ ppdiblc1 = 3.067627634691839E-13 pdiblc2 = 0.06924235339538 lpdiblc2 = -1.348171764075202E-8
+ wpdiblc2 = -3.512594260368968E-8 ppdiblc2 = 7.218006467461038E-15 pdiblcb = -0.311465201285046
+ lpdiblcb = 5.414186743199809E-10 wpdiblcb = 1.266016243394434E-7 ppdiblcb = -2.898713351652542E-16
+ drout = -0.670911346534265 ldrout = 3.475295091429687E-7 wdrout = 8.945929018259426E-7
+ pdrout = -1.860645884649742E-13 pscbe1 = 7.451439241051142E8 lpscbe1 = 11.409405513225517
+ wpscbe1 = 29.369515156729904 ppscbe1 = -6.108506718417939E-6 pscbe2 = 1.668749840172835E-7
+ lpscbe2 = -2.730318774420894E-14 wpscbe2 = -8.430990158260547E-14 ppscbe2 = 1.461791375338506E-20
+ pvag = 0 delta = 0.01 fprout = 0
+ pdits = 0 pditsl = 0 pditsd = 0
+ lambda = 0 vtl = 0 lc = 5E-9
+ xn = 3 alpha0 = 1E-10 alpha1 = 1E-10
+ beta0 = 12.3380115033282 lbeta0 = -1.351653934078148E-6 wbeta0 = -2.450913971186632E-6
+ pbeta0 = 7.236649734047544E-13 aigbacc = 0.43 bigbacc = 0.054
+ cigbacc = 0.075 nigbacc = 1 aigbinv = 0.35
+ bigbinv = 0.03 cigbinv = 6E-3 eigbinv = 1.1
+ nigbinv = 3 aigc = 0.43 bigc = 0.054
+ cigc = 0.075 aigsd = 0.43 bigsd = 0.054
+ cigsd = 0.075 dlcig = 0 nigc = 1
+ poxedge = 1 pigcd = 1 ntox = 1
+ toxref = 4.23E-9 agidl = -5.89222603784416E-8 lagidl = 1.055800817495218E-14
+ wagidl = 3.235685692646298E-14 pagidl = -5.652675224405634E-21 bgidl = 1E9
+ cgidl = 300 egidl = 0.1 noia = 1.5E42
+ noib = 0 noic = 0 em = 4.1E7
+ af = 1 ef = 1 kf = 0
+ lintnoi = -2E-7 tnoia = 2.5E7 tnoib = 0
+ ntnoi = 1 rnoia = 0.69 rnoib = 0.34
+ xpart = 0 cgso = {5.248925E-11/sw_func_tox_lv_ratio} cgdo = {5.248925E-11/sw_func_tox_lv_ratio}
+ cgbo = {0/sw_func_tox_lv_ratio} ckappas = 0.6 cf = 1.2E-11
+ clc = 1E-7 cle = 0.6 dlc = -3E-9
+ dwc = 0 vfbcv = -0.14469 noff = 3.9
+ voffcv = -0.10701 acde = 0.8 moin = 18.13
+ cgsl = {9.548271750000001E-12/sw_func_tox_lv_ratio} cgdl = {9.548271750000001E-12/sw_func_tox_lv_ratio} ijthsrev = 0.1
+ ijthsfwd = 0.1 xjbvs = 1 bvs = 12.69
+ jss = 2.1483E-5 jsws = 8.040000000000001E-10 cjs = {sw_psd_nw_cj}
+ mjs = 0.34629 mjsws = 0.29781 cjsws = {9.888891999999999E-11*sw_func_psd_nw_cj}
+ cjswgs = {2.39155046E-10*sw_func_psd_nw_cj} mjswgs = 0.9274 pbs = 0.6587
+ pbsws = 0.7418 pbswgs = 1.4338 xrcrg1 = 12
+ xrcrg2 = 1 rbpb = 50 rbpd = 50
+ rbps = 50 rbdb = 50 rbsb = 50
+ gbmin = 1E-12 tnom = 30 ute = -0.143066025781538
+ lute = 1.154412545731235E-7 wute = 7.659643428843436E-8 pute = -6.180634725666467E-14
+ kt1 = -0.704020798415384 wkt1 = 3.300735659536919E-8 kt1l = 0
+ kt2 = -0.12 ua1 = -5.445875142630204E-10 lua1 = 1.354125916142738E-16
+ wua1 = 3.725138540718098E-16 pua1 = -7.249884533206762E-23 ub1 = 3.7264E-19
+ uc1 = 2.786693462483196E-10 luc1 = -5.264121208534432E-17 wuc1 = -1.360138968276496E-16
+ puc1 = 2.818369434903908E-23 at = -6.264159844354673E5 lat = 0.118792898997563
+ wat = 0.366781661513071 pat = -6.360079153868316E-8 prt = 0
+ njs = 1.3632 xtis = 5.2 tpb = 2.0386E-3
+ tpbsw = 1.246E-3 tpbswg = 0 tcj = 1.2407E-3
+ tcjsw = 3.7357E-4 tcjswg = 2E-12 tvoff = 0
+ tvfbsdoff = 0 saref = 1.1E-6 sbref = 1.1E-6
+ wlod = 0 ku0 = 4.5E-8 kvsat = 0.5
+ kvth0 = 3.29E-8 tku0 = 0 llodku0 = 0
+ wlodku0 = 1 llodvth = 0 wlodvth = 1
+ lku0 = 0 wku0 = 2.5E-7 pku0 = 0
+ lkvth0 = 0 wkvth0 = 2E-7 pkvth0 = 0
+ stk2 = 0 lodk2 = 1 steta0 = 0
+ lodeta0 = 1

.ends sky130_fd_pr__pfet_01v8
