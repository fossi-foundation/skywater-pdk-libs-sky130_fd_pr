* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

******************************************************************
******************************************************************
*  *****************************************************
*  03/08/2021 Usman Suriono
*      Why     : New infrastructure of the ESD sky130_fd_pr__nfet_01v8 5V model.
*      What    : Converted from nhvesd model into a continuous model.
*
*  *****************************************************
*
*  ESD Nmos 5V Model
*  -----------------------------------------------------

.subckt  sky130_fd_pr__esd_nfet_g5v0d10v5 d g s b mult=1
+ 
.param  l = 1 w = 1 nf = 1 ad = 0 as = 0 pd = 0 ps = 0 nrd = {0.14/w} nrs = {0.14/w} sa = 0 sb = 0 sd = 0
+ swx_nrds = {89.1*nf/w+443.5}
* Corners and MC
+ swx_vth = {sw_vth0_sky130_fd_pr__nfet_g5v0d10v5+sw_mm_vth0_sky130_fd_pr__nfet_g5v0d10v5*mismatch_factor*MC_MM_SWITCH*AGAUSS(0,1.0,1)/sqrt(l*w*mult)+sw_vth0_sky130_fd_pr__nfet_g5v0d10v5_mc}
* legacy fitting parameters from Cypress
+ sky130_fd_pr__esd_nfet_g5v0d10v5_nfactor_diff_2 = 0.23391
+ sky130_fd_pr__esd_nfet_g5v0d10v5_k2_diff_2 = 0.010304
+ sky130_fd_pr__esd_nfet_g5v0d10v5_u0_diff_2 = 0.0012741
+ sky130_fd_pr__esd_nfet_g5v0d10v5_vth0_diff_2 = 0.013326
+ sky130_fd_pr__esd_nfet_g5v0d10v5_vsat_diff_2 = -43.451
+ sky130_fd_pr__esd_nfet_g5v0d10v5_ub_diff_2 = 3.291e-19
+ sky130_fd_pr__esd_nfet_g5v0d10v5_ua_diff_2 = -7.333e-12


Msky130_fd_pr__esd_nfet_g5v0d10v5 d g s b sky130_fd_pr__esd_nfet_g5v0d10v5_model l = {l} w = {w} ad = {ad} as = {as} pd = {pd} ps = {ps} nrd = {nrd} nrs = {nrs} sa = {sa} sb = {sb} sd = {sd} nf = {nf}
* + deltox = 0.3*(sw_tox_hv_corner - sw_tox_hv_nom) + sw_tox_hv_mc + sw_mm_tox_hv * mismatch_factor*MC_MM_SWITCH*AGAUSS(0,1.0,1)/sqrt(l*w*mult)
+ delvto = {-0.006+0.02*(1/l-1/0.55)+swx_vth*1.35}
* + mulvsat = 0.93 * (sw_vsat_sky130_fd_pr__nfet_g5v0d10v5**0.5) * (1 + 0.25*(1/l - 1/0.55))




.model sky130_fd_pr__esd_nfet_g5v0d10v5_model.0 nmos
+ 
*
* DC IV MOS PARAMETERS
*
+ lmin = 5.45e-07 lmax = 1.05e-06 wmin = 17.495e-06 wmax = 1.05e-04
+ level = 54
+ tnom = 30
+ version = 4.5
+ toxm = 1.16e-008
+ xj = 1.5e-007
+ lln = 1
+ lwn = 1
+ wln = 1
+ wwn = 1
+ lint = {3.6e-008-sw_polycd}
+ ll = 0
+ lw = 0
+ lwl = 0
+ wint = {-5.8413e-010+sw_activecd}
+ wl = 0
+ ww = 0
+ wwl = 0
+ xl = 0
+ xw = 0
+ mobmod = 0
+ binunit = 2
+ dwg = 0
+ dwb = 3.3727471e-012
* NEW BSIM4 Parameters(Model Selectors)
+ igcmod = 0
+ igbmod = 0
+ rgatemod = 0
+ rbodymod = 1
+ trnqsmod = 0
+ acnqsmod = 0
+ fnoimod = 1
+ tnoimod = 1
+ permod = 1
+ geomod = 0
+ rdsmod = 0
+ tempmod = 0
* ******
* NEW BSIM4 Parameters(4.4 Version)
+ lintnoi = 0.0
+ vfbsdoff = 0
+ lambda = 0
+ vtl = 0
+ lc = 5e-009
+ xn = 3
+ rnoia = 0.577
+ rnoib = 0.5164
+ tnoia = 1.5
+ tnoib = 3.5
* NEW BSIM4 Parameters(Process Parameters)
+ epsrox = 3.9
+ toxe = 1.16e-008
+ dtox = 0
+ ndep = 1.7e+017
+ nsd = 1e+020
+ rshg = 0.1
* ***
+ rsh = {swx_nrds}
*
*  THRESHOLD VOLTAGE PARAMETERS
*
+ vth0 = {0.814+sky130_fd_pr__esd_nfet_g5v0d10v5_vth0_diff_2}
+ k1 = 0.76281
+ k2 = {-0.081731+sky130_fd_pr__esd_nfet_g5v0d10v5_k2_diff_2}
+ k3 = 0
+ dvt0 = 0
+ dvt1 = 0.5
+ dvt2 = -0.001152
+ dvt0w = 0
+ dvt1w = 5215200
+ dvt2w = -0.036016
+ w0 = 0
+ k3b = 0
* NEW BSIM4 Parameters for Level 54
+ phin = 0
+ lpe0 = 0
+ lpeb = 0
+ vbm = -3
+ dvtp0 = 0
+ dvtp1 = 0
*
*  MOBILITY PARAMETERS
*
+ vsat = {107440+sky130_fd_pr__esd_nfet_g5v0d10v5_vsat_diff_2}
+ ua = {1.3637e-009+sky130_fd_pr__esd_nfet_g5v0d10v5_ua_diff_2}
+ ub = {1.4129e-018+sky130_fd_pr__esd_nfet_g5v0d10v5_ub_diff_2}
+ uc = 4.4957e-011
+ rdsw = 566.95
+ prwb = 0.015804
+ prwg = 5.4e-013
+ wr = 1
+ u0 = {0.066871+sky130_fd_pr__esd_nfet_g5v0d10v5_u0_diff_2}
+ a0 = 0.1054
+ keta = -0.057372
+ a1 = 0
+ a2 = 0.65972622
+ ags = 0.48
+ b0 = 0
+ b1 = 0
* NEW BSIM4 Parameters(Mobility Parameters)
+ eu = 1.67
+ rdswmin = 0
+ rdw = 0
+ rdwmin = 0
+ rsw = 0
+ rswmin = 0
* ****
*
*  SUBTHRESHOLD CURRENT PARAMETERS
*
+ voff = 0
+ nfactor = {0.114+sky130_fd_pr__esd_nfet_g5v0d10v5_nfactor_diff_2}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0
+ cit = -0.0007128
+ cdsc = 0
+ cdscb = 0
+ cdscd = 4e-012
+ eta0 = 0.21835
+ etab = -0.0031079
+ dsub = 0.5
* NEW BSIM4 Parameters(Sub-threshold parameters)
+ voffl = -4.2579486e-007
+ minv = 0
* ****
*
*  ROUT PARAMETERS
*
+ pclm = 0.23915
+ pdiblc1 = 0.09332
+ pdiblc2 = 0
+ pdiblcb = -0.26831
+ drout = 0.2822
+ pscbe1 = 5.088e+008
+ pscbe2 = 2e-008
+ pvag = 1.9901676
+ delta = 0.0445
+ alpha0 = 2.6845e-005
+ alpha1 = 0.37039
+ beta0 = 39.827
* NEW BSIM4 Parameters(ROUT Parameters)
+ fprout = 10.125
+ pdits = 0
+ pditsl = 0
+ pditsd = 0
* ***
* NEW BSIM4 Parameters(GATE INDUCED DRAIN LEAKAGE MODEL PARAMTERS)
+ agidl = 5.4829e-007
+ bgidl = 2.4214e+009
+ cgidl = 10120
+ egidl = 0.8
* ***
* NEW BSIM4 Parameters(Gate Leakage Current Parameters)
+ aigbacc = 1
+ bigbacc = 0
+ cigbacc = 0
+ nigbacc = 1
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0
+ poxedge = 1
+ pigcd = 1
+ ntox = 1
+ toxref = 1.16e-008
* ****
*
*  TEMPERATURE EFFECTS PARAMETERS
*
+ kt1 = -0.34313
+ kt2 = -0.015814
+ at = 38574
+ ute = -1.4571
+ ua1 = 3.4582e-009
+ ub1 = -3.4538e-018
+ uc1 = 4.7889e-011
+ kt1l = 0
+ prt = 0
* NEW BSIM4 Parameters(HIGH SPEED RF MODEL PARAMETERS)
+ xrcrg1 = 12
+ xrcrg2 = 1
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ rbdb = 50
+ rbsb = 50
+ gbmin = 1e-012
* ***
* NEW BSIM4 Parameters(FLICKER and THERMAL NOISE PARAMETERS)
+ noia = 2.6e+41
+ noib = 0.0
+ noic = 0.0
+ em = 4.1000000E+07
+ af = 1
+ ef = 0.89
+ kf = 0
+ ntnoi = 1
* ****
* NEW BSIM4 Parameters(LAYOUT DEPENDENT PARASITIC MODEL PARAMETERS)
+ dmcg = 0
+ dmcgt = 0
+ dmdg = 0
+ xgw = 0
+ xgl = 0
+ ngcon = 1
* ***
*
* DIODE DC IV PARAMTERS
*
* NEW BSIM4 Parameters(DIODE DC IV parameters)
+ diomod = 1
+ njs = 1.0773
+ jss = 0.000375
+ jsws = 5.84e-11
+ xtis = 2
+ bvs = 12.636
+ xjbvs = 1
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
*
*  DIODE and FET CAPACITANCE PARAMETERS
*
+ tpb = 0.001344
+ tpbsw = 0.00099005
+ tpbswg = 0
+ tcj = 0.00067434
+ tcjsw = 0.0002493
+ tcjswg = 0
+ cgdo = {3.0674e-010/sw_func_tox_hv_ratio}
+ cgso = {3.0674e-010/sw_func_tox_hv_ratio}
+ cgbo = 0
+ capmod = 2
+ xpart = 0
+ cgsl = {5e-011/sw_func_tox_hv_ratio}
+ cgdl = {5e-011/sw_func_tox_hv_ratio}
+ cf = 0
+ clc = 1e-007
+ cle = 0.6
+ dlc = {6.5995e-008-sw_polycd}
+ dwc = {sw_activecd}
+ vfbcv = -1
+ acde = 0.4176
+ moin = 15
+ noff = 4
+ voffcv = -0.4104
+ ngate = 1e+023
+ lwc = 0
+ llc = 0
+ lwlc = 0
+ wlc = 0
+ wwc = 0
+ wwlc = 0
* NEW BSIM4 Parameters(FET and DIODE capacitance parameters)
+ ckappas = 0.6
+ cjs = {0.0008512*sw_func_nsd_pw_cj}
+ mjs = 0.295
+ pbs = 0.72468
+ cjsws = {8.5204e-011*sw_func_nsd_pw_cj}
+ mjsws = 0.037586
+ pbsws = 0.29067
+ cjswgs = {5.4e-011*sw_func_nsd_pw_cj}
+ mjswgs = 0.78692
+ pbswgs = 0.54958
* *****

.ends sky130_fd_pr__esd_nfet_g5v0d10v5
