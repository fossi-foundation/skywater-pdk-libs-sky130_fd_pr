* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

*  -----------------------------------------------------
*       Base Pmos VHV DE Model
*  -----------------------------------------------------

.subckt  sky130_fd_pr__pfet_g5v0d16v0_base  d g s b  mult=1
+ l=1 w=1 
.param  nf = 1 ad = 0 as = 0 pd = 0 ps = 0 nrd = 0 nrs = 0 sa = 0 sb = 0 sd = 0

Msky130_fd_pr__pfet_g5v0d16v0_base  d g s b pvhv_model_base l = {l} w = {w} ad = {ad} as = {as} pd = {pd} ps = {ps} nrd = {nrd} nrs = {nrs*sw_rdp/sw_pw_rs} sa = {sa} sb = {sb} sd = {sd} nf = {nf}
* + deltox  = 0.3*(sw_tox_hv_corner - sw_tox_hv_nom) + sw_tox_hv_mc + sw_mm_tox_hv * mismatch_factor*MC_MM_SWITCH*AGAUSS(0,1.0,1)/sqrt(l*w*mult)
* + mulu0   = 0.95*sw_u0_sky130_fd_pr__pfet_g5v0d16v0**(-0.2*0.66/l+1.2)
+ delvto = {-0.0005+sw_vth0_sky130_fd_pr__pfet_g5v0d16v0*(0.008*2.2/l+0.992)*(0.0007*44/(w*l)+0.9993)+sw_mm_vth0_sky130_fd_pr__pfet_g5v0d16v0*mismatch_factor*MC_MM_SWITCH*AGAUSS(0,1.0,1)/sqrt(l*w*mult)+sw_vth0_sky130_fd_pr__pfet_g5v0d16v0_mc}
* + delk1   = -0.25*(sw_vth0_sky130_fd_pr__pfet_g5v0d16v0 + sw_vth0_sky130_fd_pr__pfet_g5v0d16v0_mc)
* + mulvsat = sw_vsat_sky130_fd_pr__pfet_g5v0d16v0**(-0.3*0.66/l + 1.3)




.model pvhv_model_base.1 pmos
+ level = 54 lmin = 2.16E-6 lmax = 2.02E-5 wmin = 5E-6
+ wmax = 1.01E-3 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 1 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ permod = 1 geomod = 0 rgatemod = 0
+ epsrox = 3.9 toxe = 1.16E-8 toxm = 1.16E-8
+ xj = 1.5E-7 ndep = 1.7E17 ngate = 1E23
+ nsd = 1E20 rsh = {sw_pw_rs} rshg = 0.1
+ phin = 0 wint = {0+sw_activecd} wl = 0
+ wln = 1 ww = 0 wwn = 1
+ wwl = 0 lint = {3.4453E-8-sw_polycd} ll = 0
+ lln = 1 lw = 0 lwn = 1
+ lwl = 0 llc = 0 lwc = 0
+ lwlc = 0 wlc = 0 wwc = 0
+ wwlc = 0 dwg = 0 dwb = 0
+ xl = 0 xw = 0 dmcg = 0
+ dmdg = 0 dmcgt = 0 xgw = 0
+ xgl = 0 ngcon = 1 vth0 = -1.102088
+ k1 = 0.6831 k2 = -1.3032E-3 k3 = 0
+ k3b = 0 w0 = 0 lpe0 = 1.4E-7
+ lpeb = -6.5E-8 vbm = -3 dvtp0 = 0
+ dvtp1 = 0 dvt0 = 0 dvt1 = 0.53
+ dvt2 = -0.032 dvt0w = 0 dvt1w = 5.3E6
+ dvt2w = -0.032 u0 = 2.61536E-2 ua = 2.5856E-9
+ ub = 4.5958E-19 uc = -1.22E-10 eu = 1.67
+ vsat = 7.6608E4 a0 = 0.382 ags = 0.12912
+ b0 = 4E-12 b1 = 0 keta = -0.033218
+ a1 = 0 a2 = 0.72 rdsw = 331.02
+ rdswmin = 0 rdw = 10 rdwmin = 0
+ rsw = 100 rswmin = 0 prwb = -4E-4
+ prwg = 0 wr = 1 voff = -0.1372
+ voffl = 0 minv = 0 nfactor = 0.71
+ eta0 = 0.087298 etab = -0.05 dsub = 0.3416
+ cit = 0 cdsc = 2.52E-4 cdscb = 0
+ cdscd = 0 pclm = 0.1 pdiblc1 = 0.39
+ pdiblc2 = 8.6E-3 pdiblcb = -5.4E-5 drout = 0.56
+ pscbe1 = 5.088E8 pscbe2 = 6.9452E-9 pvag = 0.504
+ delta = 8.9E-3 fprout = 0 pdits = 0
+ pditsl = 0 pditsd = 0 alpha0 = 2E-7
+ alpha1 = 1.001 beta0 = 100 aigbacc = 0.43
+ bigbacc = 0.054 cigbacc = 0.075 nigbacc = 1
+ aigbinv = 0.35 bigbinv = 0.03 cigbinv = 6E-3
+ eigbinv = 1.1 nigbinv = 3 aigc = 0.43
+ bigc = 0.054 cigc = 0.075 aigsd = 0.43
+ bigsd = 0.054 cigsd = 0.075 nigc = 1
+ poxedge = 1 pigcd = 1 ntox = 1
+ toxref = 1.16E-8 agidl = 1.65E-10 bgidl = 5.9993E9
+ cgidl = 1.394 egidl = 0.0492 noia = 6.25E41
+ noib = 3.125E26 noic = 8.75E9 em = 4.1E7
+ ef = 1 xpart = 0 cgso = {1.9771E-10/sw_func_tox_hv_ratio}
+ cgdo = {1.9771E-10/sw_func_tox_hv_ratio} cgbo = {0/sw_func_tox_hv_ratio} ckappas = 0.6
+ ckappad = 0.6 cf = 0 clc = 6.324E-9
+ cle = 0.891 dlc = -9.6826E-8 dwc = 0
+ vfbcv = -1 noff = 1.045 voffcv = -0.18151
+ acde = 0.91298 moin = 15.562 cgsl = {1.152E-12/sw_func_tox_hv_ratio}
+ cgdl = {1.1172E-12/sw_func_tox_hv_ratio} ijthsrev = 0.1 ijthsfwd = 0.1
+ xjbvs = 1 bvs = 12.69 jss = 2.1483E-5
+ jsws = 4.02E-12 jtssws = 0 cjs = {8.310E-04*sw_func_nsd_pw_cj}
+ mjs = 0.33956 mjsws = 0.24676 cjsws = {9.960545E-11*sw_func_nsd_pw_cj}
+ cjswgs = {1.47314E-10*sw_func_nsd_pw_cj} mjswgs = 0.81 pbs = 0.6587
+ pbsws = 1 pbswgs = 3 tnom = 30
+ ute = -1.6462 kt1 = -0.49308 kt1l = 1E-11
+ kt2 = 5.6338E-4 ua1 = 1.2181E-9 ub1 = -1.2412E-18
+ uc1 = 8.272E-12 at = -6.4E4 prt = 0
+ njs = 1.3632 njd = 1.0791 xtis = 10
+ xtid = 3 tpb = 1.671E-3 tpbsw = 0
+ tpbswg = 0 tcj = 9.6E-4 tcjsw = 3E-5
+ tcjswg = 0 tvoff = 0.015 saref = 2.8E-7
+ sbref = 1.19E-6 wlod = 0 ku0 = 2.218E-7
+ kvsat = 0.4 kvth0 = 5.2302E-9 tku0 = 0
+ llodku0 = 1 wlodku0 = 1 llodvth = 1
+ wlodvth = 1 lku0 = 8.7129E-7 wku0 = 0
+ pku0 = 0 lkvth0 = -4.8631E-7 wkvth0 = 5.398E-7
+ pkvth0 = 0 stk2 = 0 lodk2 = 1
+ steta0 = 0 lodeta0 = 1

.model pvhv_model_base.2 pmos
+ level = 54 lmin = 6.6E-7 lmax = 2.16E-6 wmin = 5E-6
+ wmax = 1.01E-3 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 1 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ permod = 1 geomod = 0 rgatemod = 0
+ epsrox = 3.9 toxe = 1.16E-8 toxm = 1.16E-8
+ xj = 1.5E-7 ndep = 1.7E17 ngate = 1E23
+ nsd = 1E20 rsh = {sw_pw_rs} rshg = 0.1
+ phin = 0 wint = {0+sw_activecd} wl = 0
+ wln = 1 ww = 0 wwn = 1
+ wwl = 0 lint = {3.4453E-8-sw_polycd} ll = 0
+ lln = 1 lw = 0 lwn = 1
+ lwl = 0 llc = 0 lwc = 0
+ lwlc = 0 wlc = 0 wwc = 0
+ wwlc = 0 dwg = 0 dwb = 0
+ xl = 0 xw = 0 dmcg = 0
+ dmdg = 0 dmcgt = 0 xgw = 0
+ xgl = 0 ngcon = 1 vth0 = -1.112786
+ lvth0 = 2.237055E-8 k1 = 0.6831 k2 = -1.3032E-3
+ k3 = 0 k3b = 0 w0 = 0
+ lpe0 = 1.4E-7 lpeb = -6.5E-8 vbm = -3
+ dvtp0 = 0 dvtp1 = 0 dvt0 = 0
+ dvt1 = 0.53 dvt2 = -0.032 dvt0w = 0
+ dvt1w = 5.3E6 dvt2w = -0.032 u0 = 2.68468E-2
+ lu0 = -1.449455E-9 ua = 2.5856E-9 ub = 4.5958E-19
+ uc = -1.22E-10 eu = 1.67 vsat = 7.6608E4
+ a0 = 0.382 ags = 0.12912 b0 = 4E-12
+ b1 = 0 keta = -0.033218 a1 = 0
+ a2 = 0.72 rdsw = 331.02 rdswmin = 0
+ rdw = 10 rdwmin = 0 rsw = 100
+ rswmin = 0 prwb = -4E-4 prwg = 0
+ wr = 1 voff = -0.1372 voffl = 0
+ minv = 0 nfactor = 0.71 eta0 = 0.087298
+ etab = -0.05 dsub = 0.3416 cit = 0
+ cdsc = 2.52E-4 cdscb = 0 cdscd = 0
+ pclm = 0.1 pdiblc1 = 0.39 pdiblc2 = 8.6E-3
+ pdiblcb = -5.4E-5 drout = 0.56 pscbe1 = 5.088E8
+ pscbe2 = 6.9452E-9 pvag = 0.504 delta = 8.9E-3
+ fprout = 0 pdits = 0 pditsl = 0
+ pditsd = 0 alpha0 = 2E-7 alpha1 = 1.001
+ beta0 = 100 aigbacc = 0.43 bigbacc = 0.054
+ cigbacc = 0.075 nigbacc = 1 aigbinv = 0.35
+ bigbinv = 0.03 cigbinv = 6E-3 eigbinv = 1.1
+ nigbinv = 3 aigc = 0.43 bigc = 0.054
+ cigc = 0.075 aigsd = 0.43 bigsd = 0.054
+ cigsd = 0.075 nigc = 1 poxedge = 1
+ pigcd = 1 ntox = 1 toxref = 1.16E-8
+ agidl = 1.65E-10 bgidl = 5.9993E9 cgidl = 1.394
+ egidl = 0.0492 noia = 6.25E41 noib = 3.125E26
+ noic = 8.75E9 em = 4.1E7 ef = 1
+ xpart = 0 cgso = {1.9771E-10/sw_func_tox_hv_ratio} cgdo = {1.9771E-10/sw_func_tox_hv_ratio}
+ cgbo = {0/sw_func_tox_hv_ratio} ckappas = 0.6 ckappad = 0.6
+ cf = 0 clc = 6.324E-9 cle = 0.891
+ dlc = -9.6826E-8 dwc = 0 vfbcv = -1
+ noff = 1.045 voffcv = -0.18151 acde = 0.91298
+ moin = 15.562 cgsl = {1.152E-12/sw_func_tox_hv_ratio} cgdl = {1.1172E-12/sw_func_tox_hv_ratio}
+ ijthsrev = 0.1 ijthsfwd = 0.1 xjbvs = 1
+ bvs = 12.69 jss = 2.1483E-5 jsws = 4.02E-12
+ jtssws = 0 cjs = {8.310E-04*sw_func_nsd_pw_cj} mjs = 0.33956
+ mjsws = 0.24676 cjsws = {9.960545E-11*sw_func_nsd_pw_cj} cjswgs = {1.47314E-10*sw_func_nsd_pw_cj}
+ mjswgs = 0.81 pbs = 0.6587 pbsws = 1
+ pbswgs = 3 tnom = 30 ute = -1.6462
+ kt1 = -0.49308 kt1l = 1E-11 kt2 = 5.6338E-4
+ ua1 = 1.2181E-9 ub1 = -1.2412E-18 uc1 = 8.272E-12
+ at = -6.4E4 prt = 0 njs = 1.3632
+ njd = 1.0791 xtis = 10 xtid = 3
+ tpb = 1.671E-3 tpbsw = 0 tpbswg = 0
+ tcj = 9.6E-4 tcjsw = 3E-5 tcjswg = 0
+ tvoff = 0.015 saref = 2.8E-7 sbref = 1.19E-6
+ wlod = 0 ku0 = 2.218E-7 kvsat = 0.4
+ kvth0 = 5.2302E-9 tku0 = 0 llodku0 = 1
+ wlodku0 = 1 llodvth = 1 wlodvth = 1
+ lku0 = 8.7129E-7 wku0 = 0 pku0 = 0
+ lkvth0 = -4.8631E-7 wkvth0 = 5.398E-7 pkvth0 = 0
+ stk2 = 0 lodk2 = 1 steta0 = 0
+ lodeta0 = 1

.ends sky130_fd_pr__pfet_g5v0d16v0_base
