* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

******************************************************************
******************************************************************
*  *****************************************************
*  05/04/2021 Usman Suriono
*      Why     : To follow sky130_fd_pr__nfet_05v0_nvt process monte carlo
*      What    : Adjusted the VTH monte carlo parameter.
*  04/22/2021 Usman Suriono
*      Why     : New infrastructure of the ESD sky130_fd_pr__nfet_01v8 native 5V model.
*      What    : Converted from nhvnativeesd model into a continuous model.
*                Replaced rsh from 1 to calculated rsh from the original model.
*                PDK netlist nrd/nrs = ratio of distance the middle of the contact to Gate.
*                Changed the parasitic diode from internal dimension calculation
*                to receive it from PDK
*
*  *****************************************************
*
*  ESD Nmos Native 5V Model
*  -----------------------------------------------------

.subckt  sky130_fd_pr__esd_nfet_05v0_nvt d g s b mult=1
+ 
.param  l = 1 w = 1 nf = 1 ad = 0 as = 0 pd = 0 ps = 0 nrd = {0.14/w} nrs = {0.14/w} sa = 0 sb = 0 sd = 0
+ swx_nrds = {89.1*nf/w+443.5}
*   Legacy parameter fitting from Cypress
+ sky130_fd_pr__nfet_05v0_nvt_dlc_diff = -1.5781e-08
+ sky130_fd_pr__nfet_05v0_nvt_ub_diff_2 = -1.5224e-18
+ sky130_fd_pr__nfet_05v0_nvt_nfactor_diff_2 = -0.044586
+ sky130_fd_pr__nfet_05v0_nvt_k2_diff_2 = 0.0015915
+ sky130_fd_pr__nfet_05v0_nvt_u0_diff_2 = -0.008363
+ sky130_fd_pr__nfet_05v0_nvt_ua_diff_2 = -3.3419e-11
+ sky130_fd_pr__nfet_05v0_nvt_vsat_diff_2 = -2848.5
+ sky130_fd_pr__nfet_05v0_nvt_vth0_diff_2 = -0.0011931
** NHVNATIVE NMOS STRESS PARAMS ***
+ sky130_fd_pr__nfet_05v0_nvt_wkvth0_diff = 0.8e-6
+ sky130_fd_pr__nfet_05v0_nvt_kvth0_diff = -7e-9
+ sky130_fd_pr__nfet_05v0_nvt_ku0_diff = -3e-8
+ sky130_fd_pr__nfet_05v0_nvt_wku0_diff = 0.2e-6
+ sky130_fd_pr__nfet_05v0_nvt_kvsat_diff = 0.4



Msky130_fd_pr__esd_nfet_05v0_nvt d g s b sky130_fd_pr__esd_nfet_05v0_nvt_model l = {l} w = {w} ad = {ad} as = {as} pd = {pd} ps = {ps} nrd = {nrd} nrs = {nrs} sa = {sa} sb = {sb} sd = {sd} nf = {nf}
* + deltox = 0.3*(sw_tox_hv_corner - sw_tox_hv_nom) + sw_tox_hv_mc + sw_mm_tox_hv * mismatch_factor*MC_MM_SWITCH*AGAUSS(0,1.0,1)/sqrt(l*w*mult)
+ delvto = {sw_vth0_sky130_fd_pr__nfet_01v8_nat+sw_mm_vth0_sky130_fd_pr__nfet_01v8_nat*mismatch_factor*MC_MM_SWITCH*AGAUSS(0,1.0,1)/sqrt(l*w*mult)+sw_vth0_sky130_fd_pr__nfet_01v8_nat_mc*3}
* + mulu0  = sw_u0_sky130_fd_pr__nfet_01v8_nat



.model sky130_fd_pr__esd_nfet_05v0_nvt_model nmos 
*
* DC IV MOS PARAMETERS
*
+ lmin = 8.95e-07 lmax = 4.05e-06 wmin = 9.995e-06 wmax = 1.0005e-03
+ level = 54
+ tnom = 30
+ version = 4.5
+ toxm = 1.16e-008
+ xj = 1.5e-007
+ lln = 1
+ lwn = 1
+ wln = 1
+ wwn = 1
+ lint = {6.93e-008-sw_polycd}
+ ll = 0
+ lw = 0
+ lwl = 0
+ wint = {4.5e-008+sw_activecd}
+ wl = 0
+ ww = 0
+ wwl = 0
+ xl = 0
+ xw = 0
+ mobmod = 0
+ binunit = 2
+ dwg = -4.6e-009
+ dwb = 1.92e-009
* NEW BSIM4 Parameters(Model Selectors)
+ igcmod = 0
+ igbmod = 0
+ rgatemod = 0
+ rbodymod = 1
+ trnqsmod = 0
+ acnqsmod = 0
+ fnoimod = 1
+ tnoimod = 1
+ permod = 1
+ geomod = 0
+ rdsmod = 0
+ tempmod = 0
* ******
* NEW BSIM4 Parameters(4.4 Version)
+ lintnoi = 0.0
+ vfbsdoff = 0
+ lambda = 0
+ vtl = 0
+ lc = 5e-009
+ xn = 3
+ rnoia = 0.8
+ rnoib = 0.38
+ tnoia = 7.6e6
+ tnoib = 7.2e6
* NEW BSIM4 Parameters(Process Parameters)
+ epsrox = 3.9
+ toxe = 1.16e-008
+ dtox = 0
+ ndep = 1.7e+017
+ nsd = 1e+020
+ rshg = 0.1
* ***
+ rsh = {swx_nrds}
*
*  THRESHOLD VOLTAGE PARAMETERS
*
+ vth0 = {0.062+sky130_fd_pr__nfet_05v0_nvt_vth0_diff_2}
+ k1 = 0.364
+ k2 = {0.038817+sky130_fd_pr__nfet_05v0_nvt_k2_diff_2}
+ k3 = 1.4
+ dvt0 = 5.7
+ dvt1 = 0.21851
+ dvt2 = 0.04
+ dvt0w = 7.7
+ dvt1w = 1272000
+ dvt2w = -0.032
+ w0 = 0
+ k3b = -0.58
* NEW BSIM4 Parameters for Level 54
+ phin = 0
+ lpe0 = -1.2362266e-014
+ lpeb = 0
+ vbm = -3
+ dvtp0 = 0
+ dvtp1 = 0
*
*  MOBILITY PARAMETERS
*
+ vsat = {74500+sky130_fd_pr__nfet_05v0_nvt_vsat_diff_2}
+ ua = {9.1406e-010+sky130_fd_pr__nfet_05v0_nvt_ua_diff_2}
+ ub = {1.2863e-018+sky130_fd_pr__nfet_05v0_nvt_ub_diff_2}
+ uc = 3.2583e-011
+ rdsw = 430
+ prwb = 0
+ prwg = 1e-012
+ wr = 1
+ u0 = {0.050801+sky130_fd_pr__nfet_05v0_nvt_u0_diff_2}
+ a0 = 0.08
+ keta = -0.019904
+ a1 = 0
+ a2 = 0.96293372
+ ags = 0.87995
+ b0 = 3.3993e-007
+ b1 = 0
* NEW BSIM4 Parameters(Mobility Parameters)
+ eu = 1.67
+ rdswmin = 0
+ rdw = 0
+ rdwmin = 0
+ rsw = 0
+ rswmin = 0
* ****
*
*  SUBTHRESHOLD CURRENT PARAMETERS
*
+ voff = 0
+ nfactor = {0.63313+sky130_fd_pr__nfet_05v0_nvt_nfactor_diff_2}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0
+ cit = 9.2584123e-008
+ cdsc = 0
+ cdscb = 1.4150948e-007
+ cdscd = 1.5e-005
+ eta0 = 9
+ etab = -0.00021692
+ dsub = 0.42
* NEW BSIM4 Parameters(Sub-threshold parameters)
+ voffl = 1.9445332e-008
+ minv = 0
* ****
*
*  ROUT PARAMETERS
*
+ pclm = 0.11748
+ pdiblc1 = 8.833e-007
+ pdiblc2 = 0.0002
+ pdiblcb = 0
+ drout = 0.13139
+ pscbe1 = 2.4476e+008
+ pscbe2 = 3.84e-009
+ pvag = 4.5419436
+ delta = 0.007
+ alpha0 = 2.1079e-006
+ alpha1 = 0.1232
+ beta0 = 25.668
* NEW BSIM4 Parameters(ROUT Parameters)
+ fprout = 0
+ pdits = 0.0002
+ pditsl = 0
+ pditsd = 0
* ***
* NEW BSIM4 Parameters(GATE INDUCED DRAIN LEAKAGE MODEL PARAMTERS)
+ agidl = 0
+ bgidl = 2.3e+009
+ cgidl = 0.5
+ egidl = 0.8
* ***
* NEW BSIM4 Parameters(Gate Leakage Current Parameters)
+ aigbacc = 1
+ bigbacc = 0
+ cigbacc = 0
+ nigbacc = 1
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0
+ poxedge = 1
+ pigcd = 1
+ ntox = 1
+ toxref = 1.16e-008
* ****
*
*  TEMPERATURE EFFECTS PARAMETERS
*
+ kt1 = -0.37322
+ kt2 = -0.01144
+ at = 19488
+ ute = -1.464
+ ua1 = 1e-009
+ ub1 = -7.128e-019
+ uc1 = 1e-011
+ kt1l = 0
+ prt = 0
* NEW BSIM4 Parameters(HIGH SPEED RF MODEL PARAMETERS)
+ xrcrg1 = 12
+ xrcrg2 = 1
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ rbdb = 50
+ rbsb = 50
+ gbmin = 1e-012
* ***
* NEW BSIM4 Parameters(FLICKER and THERMAL NOISE PARAMETERS)
+ noia = 2.5e+41
+ noib = 0.0
+ noic = 0.0
+ em = 4.1000000E+07
+ af = 1
+ ef = 1.0
+ kf = 0
+ ntnoi = 1
* ****
* NEW BSIM4 Parameters(LAYOUT DEPENDENT PARASITIC MODEL PARAMETERS)
+ dmcg = 0
+ dmcgt = 0
+ dmdg = 0
+ xgw = 0
+ xgl = 0
+ ngcon = 1
* ***
*
* DIODE DC IV PARAMTERS
*
* NEW BSIM4 Parameters(DIODE DC IV parameters)
+ diomod = 1
+ njs = 1.5764
+ jss = 0.00042966
+ jsws = 8.040000000000001e-10
+ xtis = 0
+ bvs = 12.69
+ xjbvs = 1
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
*
*  DIODE and FET CAPACITANCE PARAMETERS
*
+ tpb = 0.0019685
+ tpbsw = 0.001
+ tpbswg = 0
+ tcj = 0.00083
+ tcjsw = 0
+ tcjswg = 0
+ cgdo = {3.473e-010/sw_func_tox_hv_ratio*7.7117e-01}
+ cgso = {3.473e-010/sw_func_tox_hv_ratio*7.7117e-01}
+ cgbo = 0
+ capmod = 2
+ xpart = 0
+ cgsl = {5e-011/sw_func_tox_hv_ratio*7.7117e-01}
+ cgdl = {5e-011/sw_func_tox_hv_ratio*7.7117e-01}
+ cf = 0
+ clc = 1e-007
+ cle = 0.6
+ dlc = {7.6493e-008+sky130_fd_pr__nfet_05v0_nvt_dlc_diff-sw_polycd}
+ dwc = {sw_activecd}
+ vfbcv = -1
+ acde = 1.16
+ moin = 15
+ noff = 4
+ voffcv = 0.216
+ ngate = 1e+023
+ lwc = 0
+ llc = 0
+ lwlc = 0
+ wlc = 0
+ wwc = 0
+ wwlc = 0
* NEW BSIM4 Parameters(FET and DIODE capacitance parameters)
+ ckappas = 0.6
+ cjs = {0.0008602*9.7602e-01*sw_func_nsd_pw_cj}
+ mjs = 0.28329
+ pbs = 0.66345
+ cjsws = {8.5152e-011*sw_func_nsd_pw_cj}
+ mjsws = 0.057926
+ pbsws = 1
+ cjswgs = {3.58e-011*sw_func_nsd_pw_cj}
+ mjswgs = 0.33
+ pbswgs = 0.2442
*
* STRESS PARAMETERS
*
+ saref = 2.54e-06
+ sbref = 2.54e-06
+ wlod = 0
+ kvth0 = {0+sky130_fd_pr__nfet_05v0_nvt_kvth0_diff}
+ lkvth0 = 0
+ wkvth0 = {0+sky130_fd_pr__nfet_05v0_nvt_wkvth0_diff}
+ pkvth0 = 0
+ llodvth = 0
+ wlodvth = 1
+ stk2 = 0
+ lodk2 = 1
+ lodeta0 = 1
+ ku0 = {0+sky130_fd_pr__nfet_05v0_nvt_ku0_diff}
+ lku0 = 0
+ wku0 = {0+sky130_fd_pr__nfet_05v0_nvt_wku0_diff}
+ pku0 = 0
+ llodku0 = 0
+ wlodku0 = 1
+ kvsat = {0+sky130_fd_pr__nfet_05v0_nvt_kvsat_diff}
+ steta0 = 0
+ tku0 = 0

.ends sky130_fd_pr__esd_nfet_05v0_nvt
* *****
