* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

******************************************************************
******************************************************************
*  *****************************************************
*  04/21/2021 Usman Suriono
*      Why     : New scalable sky130_fd_pr__nfet_01v8 low VT model
*      What    : Converted from discrete nlowvt models
*                Replaced rsh from 1 to calculated rsh from the original model.
*                PDK netlist nrd/nrs = ratio of distance the middle of the contact to Gate.
*
*  *****************************************************
*
*  Nmos Low VT Model
*  -----------------------------------------------------

.subckt  sky130_fd_pr__nfet_01v8_lvt  d g s b  mult=1
+ 
.param  l = 1 w = 1 nf = 1 ad = 0 as = 0 pd = 0 ps = 0 nrd = {0.14/w} nrs = {0.14/w} sa = 0 sb = 0 sd = 0
+ swx_nrds = {89.1*nf/w+443.5}
+ swx_vth = {sw_vth0_sky130_fd_pr__nfet_01v8_lvt+sw_vth0_sky130_fd_pr__nfet_01v8_lvt_mc}

Msky130_fd_pr__nfet_01v8_lvt  d g s b nlowvt_model l = {l} w = {w} ad = {ad} as = {as} pd = {pd} ps = {ps} nrd = {nrd} nrs = {nrs} sa = {sa} sb = {sb} sd = {sd} nf = {nf}
* + deltox = 0.3*(sw_tox_lv_corner - sw_tox_lv_nom) + sw_tox_lv_mc + sw_mm_tox_lv * mismatch_factor*MC_MM_SWITCH*AGAUSS(0,1.0,1)/sqrt(l*w*mult)
* + mulu0  = sw_u0_sky130_fd_pr__nfet_01v8_lvt
+ delvto = {swx_vth*(0.020*8/l+0.980)*(0.017*7/w+0.983)*(0.0007*56/(w*l)+0.9993)+sw_mm_vth0_sky130_fd_pr__nfet_01v8_lvt*mismatch_factor*MC_MM_SWITCH*AGAUSS(0,1.0,1)/sqrt(l*w*mult)}




.model nlowvt_model.1 nmos
+ level = 54 lmin = 8E-6 lmax = 2.02E-5 wmin = 7E-6
+ wmax = 1.01E-3 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 4.148E-9
+ toxm = 4.148E-9 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 9.999999999999999E22 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {2.6E-8+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {1.2025E-8-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = -1.33E-8 dwb = -1.08E-8 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = 0.417908 vfb = 0
+ k1 = 0.47213 k2 = -0.033282 k3 = 1.65
+ k3b = 1.6 w0 = 1E-7 lpe0 = 2.3802E-7
+ lpeb = -4.9152E-8 vbm = -3 dvtp0 = 0
+ dvtp1 = 0 dvt0 = 0.07665 dvt1 = 0.1252
+ dvt2 = -0.05637 dvt0w = 0 dvt1w = 5.3E6
+ dvt2w = -0.032 vfbsdoff = 0 u0 = 0.03198837
+ ua = -1.3015602E-9 ub = 2.67551E-18 uc = 7.0152E-11
+ ud = 0 up = 0 lp = 1
+ eu = 1.67 vsat = 1.6114E5 a0 = 1.9598449
+ ags = 0.5317926 b0 = 0 b1 = 0
+ keta = 0 a1 = 0 a2 = 0.38689047
+ rdsw = 103.65 rdswmin = 0 rdw = 0
+ rdwmin = 0 rsw = 0 rswmin = 0
+ prwb = 0 prwg = 0 wr = 1
+ voff = -0.11559919 voffl = 0 minv = 0
+ nfactor = 1.1019079 eta0 = 0.08 etab = -0.07
+ dsub = 0.56 cit = 1E-5 cdsc = 3.8556E-37
+ cdscb = -1.1484E-4 cdscd = 4.7984E-6 pclm = 0.2
+ pdiblc1 = 0.39 pdiblc2 = 4.7977E-3 pdiblcb = 0
+ drout = 3.4946 pscbe1 = 4.5E8 pscbe2 = 1E-8
+ pvag = 0 delta = 0.01 fprout = 0
+ pdits = 1.4427E-15 pditsl = 0 pditsd = 0
+ lambda = 0 vtl = 0 lc = 0
+ xn = 0 alpha0 = 8.4345657E-5 alpha1 = 0
+ beta0 = 17.822982 aigbacc = 1 bigbacc = 0
+ cigbacc = 0 nigbacc = 1 aigbinv = 0.35
+ bigbinv = 0.03 cigbinv = 6E-3 eigbinv = 1.1
+ nigbinv = 3 aigc = 0.43 bigc = 0.054
+ cigc = 0.075 aigsd = 0.43 bigsd = 0.054
+ cigsd = 0.075 dlcig = 0 nigc = 1
+ poxedge = 1 pigcd = 1 ntox = 1
+ toxref = 4.148E-9 agidl = 0 bgidl = 2.3E9
+ cgidl = 0.5 egidl = 0.8 noia = 9E41
+ noib = 1E27 noic = 8E11 em = 4.1E7
+ af = 1 ef = 1.2 kf = 0
+ lintnoi = -3E-7 tnoia = 2.5E7 tnoib = 9.9E6
+ ntnoi = 1 rnoia = 0.912 rnoib = 0.26
+ xpart = 0 cgso = {2.392894381E-10/sw_func_tox_lv_ratio} cgdo = {2.392894381E-10/sw_func_tox_lv_ratio}
+ cgbo = {1E-14/sw_func_tox_lv_ratio} ckappas = 0.6 cf = 1E-14
+ clc = 1E-7 cle = 0.6 dlc = 1.21071E-8
+ dwc = 2.6E-8 vfbcv = -1 noff = 3.8661
+ voffcv = -0.16994 acde = 0.38008 moin = 23.81
+ cgsl = {2.310725E-11/sw_func_tox_lv_ratio} cgdl = {2.310725E-11/sw_func_tox_lv_ratio} ijthsrev = 0.1
+ ijthsfwd = 0.1 xjbvs = 1 bvs = 11.9
+ jss = 2.75E-3 jsws = 6E-10 cjs = {1.210E-03*sw_func_nsd_pw_cj}
+ mjs = 0.42197 mjsws = 1E-3 cjsws = {3.230311424E-11*sw_func_nsd_pw_cj}
+ cjswgs = {1.795291232E-10*sw_func_nsd_pw_cj} mjswgs = 0.8 pbs = 0.7477
+ pbsws = 0.1 pbswgs = 0.79644 xrcrg1 = 12
+ xrcrg2 = 1 rbpb = 50 rbpd = 50
+ rbps = 50 rbdb = 50 rbsb = 50
+ gbmin = 1E-12 tnom = 30 ute = -1.0777
+ kt1 = -0.25364 kt1l = 0 kt2 = -0.034423
+ ua1 = 2.6823E-9 ub1 = -2.4433E-18 uc1 = -1.9223E-11
+ at = 3.3308E5 prt = 0 njs = 1.2928
+ xtis = 2 tpb = 1.2287E-3 tpbsw = 0
+ tpbswg = 0 tcj = 7.92E-4 tcjsw = 1E-5
+ tcjswg = 0 tvoff = 0 tvfbsdoff = 0
+ saref = 3E-6 sbref = 3E-6 wlod = 0
+ ku0 = -2.7E-8 kvsat = 0.2 kvth0 = 7.9E-9
+ tku0 = 0 llodku0 = 0 wlodku0 = 1
+ llodvth = 0 wlodvth = 1 lku0 = 0
+ wku0 = 0 pku0 = 0 lkvth0 = 0
+ wkvth0 = 3E-7 pkvth0 = 0 stk2 = 0
+ lodk2 = 1 steta0 = 0 lodeta0 = 1

.model nlowvt_model.2 nmos
+ level = 54 lmin = 4E-6 lmax = 8E-6 wmin = 7E-6
+ wmax = 1.01E-3 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 4.148E-9
+ toxm = 4.148E-9 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 9.999999999999999E22 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {2.6E-8+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {1.2025E-8-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = -1.33E-8 dwb = -1.08E-8 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = 0.417908 vfb = 0
+ k1 = 0.47213 k2 = -0.033282 k3 = 1.65
+ k3b = 1.6 w0 = 1E-7 lpe0 = 2.3802E-7
+ lpeb = -4.9152E-8 vbm = -3 dvtp0 = 0
+ dvtp1 = 0 dvt0 = 0.07665 dvt1 = 0.1252
+ dvt2 = -0.05637 dvt0w = 0 dvt1w = 5.3E6
+ dvt2w = -0.032 vfbsdoff = 0 u0 = 0.03198837
+ ua = -1.3015602E-9 ub = 2.67551E-18 uc = 7.0152E-11
+ ud = 0 up = 0 lp = 1
+ eu = 1.67 vsat = 1.6114E5 a0 = 1.9598449
+ ags = 0.5317926 b0 = 0 b1 = 0
+ keta = 0 a1 = 0 a2 = 0.38689047
+ rdsw = 103.65 rdswmin = 0 rdw = 0
+ rdwmin = 0 rsw = 0 rswmin = 0
+ prwb = 0 prwg = 0 wr = 1
+ voff = -0.11559919 voffl = 0 minv = 0
+ nfactor = 1.1019079 eta0 = 0.08 etab = -0.07
+ dsub = 0.56 cit = 1E-5 cdsc = 3.8556E-37
+ cdscb = -1.1484E-4 cdscd = 4.7984E-6 pclm = 0.2
+ pdiblc1 = 0.39 pdiblc2 = 4.7977E-3 pdiblcb = 0
+ drout = 3.4946 pscbe1 = 4.5E8 pscbe2 = 1E-8
+ pvag = 0 delta = 0.01 fprout = 0
+ pdits = 1.4427E-15 pditsl = 0 pditsd = 0
+ lambda = 0 vtl = 0 lc = 0
+ xn = 0 alpha0 = 8.4345657E-5 alpha1 = 0
+ beta0 = 17.822982 aigbacc = 1 bigbacc = 0
+ cigbacc = 0 nigbacc = 1 aigbinv = 0.35
+ bigbinv = 0.03 cigbinv = 6E-3 eigbinv = 1.1
+ nigbinv = 3 aigc = 0.43 bigc = 0.054
+ cigc = 0.075 aigsd = 0.43 bigsd = 0.054
+ cigsd = 0.075 dlcig = 0 nigc = 1
+ poxedge = 1 pigcd = 1 ntox = 1
+ toxref = 4.148E-9 agidl = 0 bgidl = 2.3E9
+ cgidl = 0.5 egidl = 0.8 noia = 9E41
+ noib = 1E27 noic = 8E11 em = 4.1E7
+ af = 1 ef = 1.2 kf = 0
+ lintnoi = -3E-7 tnoia = 2.5E7 tnoib = 9.9E6
+ ntnoi = 1 rnoia = 0.912 rnoib = 0.26
+ xpart = 0 cgso = {2.392894381E-10/sw_func_tox_lv_ratio} cgdo = {2.392894381E-10/sw_func_tox_lv_ratio}
+ cgbo = {1E-14/sw_func_tox_lv_ratio} ckappas = 0.6 cf = 1E-14
+ clc = 1E-7 cle = 0.6 dlc = 1.21071E-8
+ dwc = 2.6E-8 vfbcv = -1 noff = 3.8661
+ voffcv = -0.16994 acde = 0.38008 moin = 23.81
+ cgsl = {2.310725E-11/sw_func_tox_lv_ratio} cgdl = {2.310725E-11/sw_func_tox_lv_ratio} ijthsrev = 0.1
+ ijthsfwd = 0.1 xjbvs = 1 bvs = 11.9
+ jss = 2.75E-3 jsws = 6E-10 cjs = {1.210E-03*sw_func_nsd_pw_cj}
+ mjs = 0.42197 mjsws = 1E-3 cjsws = {3.230311424E-11*sw_func_nsd_pw_cj}
+ cjswgs = {1.795291232E-10*sw_func_nsd_pw_cj} mjswgs = 0.8 pbs = 0.7477
+ pbsws = 0.1 pbswgs = 0.79644 xrcrg1 = 12
+ xrcrg2 = 1 rbpb = 50 rbpd = 50
+ rbps = 50 rbdb = 50 rbsb = 50
+ gbmin = 1E-12 tnom = 30 ute = -1.0777
+ kt1 = -0.25364 kt1l = 0 kt2 = -0.034423
+ ua1 = 2.6823E-9 ub1 = -2.4433E-18 uc1 = -1.9223E-11
+ at = 3.3308E5 prt = 0 njs = 1.2928
+ xtis = 2 tpb = 1.2287E-3 tpbsw = 0
+ tpbswg = 0 tcj = 7.92E-4 tcjsw = 1E-5
+ tcjswg = 0 tvoff = 0 tvfbsdoff = 0
+ saref = 3E-6 sbref = 3E-6 wlod = 0
+ ku0 = -2.7E-8 kvsat = 0.2 kvth0 = 7.9E-9
+ tku0 = 0 llodku0 = 0 wlodku0 = 1
+ llodvth = 0 wlodvth = 1 lku0 = 0
+ wku0 = 0 pku0 = 0 lkvth0 = 0
+ wkvth0 = 3E-7 pkvth0 = 0 stk2 = 0
+ lodk2 = 1 steta0 = 0 lodeta0 = 1

.model nlowvt_model.3 nmos
+ level = 54 lmin = 2E-6 lmax = 4E-6 wmin = 7E-6
+ wmax = 1.01E-3 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 4.148E-9
+ toxm = 4.148E-9 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 9.999999999999999E22 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {2.6E-8+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {1.2025E-8-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = -1.33E-8 dwb = -1.08E-8 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = 0.4045856511125 lvth0 = 5.296899305925568E-8
+ vfb = 0 k1 = 0.5133680765 lk1 = -1.63960530260175E-7
+ k2 = -0.0480776172075 lk2 = 5.882663423615963E-8 k3 = 1.65
+ k3b = 1.6 w0 = 1E-7 lpe0 = 2.3802E-7
+ lpeb = -4.9152E-8 vbm = -3 dvtp0 = 0
+ dvtp1 = 0 dvt0 = 0.07665 dvt1 = 0.1252
+ dvt2 = -0.05637 dvt0w = 0 dvt1w = 5.3E6
+ dvt2w = -0.032 vfbsdoff = 0 u0 = 0.02987772936825
+ lu0 = 8.39180161980641E-9 ua = -1.37739592603125E-9 lua = 3.015190549139488E-16
+ ub = 2.6577857285E-18 lub = 7.047081727042592E-26 uc = 6.739258582500001E-11
+ luc = 1.097129278909124E-17 ud = 0 up = 0
+ lp = 1 eu = 1.67 vsat = 2.75398320775E5
+ lvsat = -0.454285370485361 a0 = 1.9486352368525 la0 = 4.45690601913023E-8
+ ags = -0.40111504464 lags = 3.709194149706409E-6 b0 = 0
+ b1 = 0 keta = 0.18231102675 lketa = -7.248595268066627E-7
+ a1 = 0 a2 = 0.38689047 rdsw = 103.65
+ rdswmin = 0 rdw = 0 rdwmin = 0
+ rsw = 0 rswmin = 0 prwb = 0
+ prwg = 0 wr = 1 voff = -0.11530539587425
+ lvoff = -1.168110754275678E-9 voffl = 0 minv = 0
+ nfactor = 0.8597940549175 lnfactor = 9.626325423557661E-7 eta0 = 0.1585440125
+ leta0 = -3.122870664993751E-7 etab = -0.1386642625 letab = 2.730056744868751E-7
+ dsub = 0.833695236578 ldsub = -1.0881985758723E-6 cit = 1E-5
+ cdsc = 3.8556E-37 cdscb = -1.1484E-4 cdscd = 4.7984E-6
+ pclm = 0.1702619525 lpclm = 1.18236989957625E-7 pdiblc1 = 0.39
+ pdiblc2 = 9.50722944999999E-4 lpdiblc2 = 1.529538842182725E-8 pdiblcb = 0
+ drout = 3.4946 pscbe1 = 4.5E8 pscbe2 = 1E-8
+ pvag = 0 delta = 0.01 fprout = 0
+ pdits = 1.4427E-15 pditsl = 0 pditsd = 0
+ lambda = 0 vtl = 0 lc = 0
+ xn = 0 alpha0 = 4.340992752532498E-5 lalpha0 = 1.627584136048341E-10
+ alpha1 = 0 beta0 = 14.391129316574998 lbeta0 = 1.364487467666363E-5
+ aigbacc = 1 bigbacc = 0 cigbacc = 0
+ nigbacc = 1 aigbinv = 0.35 bigbinv = 0.03
+ cigbinv = 6E-3 eigbinv = 1.1 nigbinv = 3
+ aigc = 0.43 bigc = 0.054 cigc = 0.075
+ aigsd = 0.43 bigsd = 0.054 cigsd = 0.075
+ dlcig = 0 nigc = 1 poxedge = 1
+ pigcd = 1 ntox = 1 toxref = 4.148E-9
+ agidl = 0 bgidl = 2.3E9 cgidl = 0.5
+ egidl = 0.8 noia = 9E41 noib = 1E27
+ noic = 8E11 em = 4.1E7 af = 1
+ ef = 1.2 kf = 0 lintnoi = -3E-7
+ tnoia = 2.5E7 tnoib = 9.9E6 ntnoi = 1
+ rnoia = 0.912 rnoib = 0.26 xpart = 0
+ cgso = {2.392894381E-10/sw_func_tox_lv_ratio} cgdo = {2.392894381E-10/sw_func_tox_lv_ratio} cgbo = {1E-14/sw_func_tox_lv_ratio}
+ ckappas = 0.6 cf = 1E-14 clc = 1E-7
+ cle = 0.6 dlc = 1.21071E-8 dwc = 2.6E-8
+ vfbcv = -1 noff = 3.8661 voffcv = -0.16994
+ acde = 0.38008 moin = 23.81 cgsl = {2.310725E-11/sw_func_tox_lv_ratio}
+ cgdl = {2.310725E-11/sw_func_tox_lv_ratio} ijthsrev = 0.1 ijthsfwd = 0.1
+ xjbvs = 1 bvs = 11.9 jss = 2.75E-3
+ jsws = 6E-10 cjs = {1.210E-03*sw_func_nsd_pw_cj} mjs = 0.42197
+ mjsws = 1E-3 cjsws = {3.230311424E-11*sw_func_nsd_pw_cj} cjswgs = {1.795291232E-10*sw_func_nsd_pw_cj}
+ mjswgs = 0.8 pbs = 0.7477 pbsws = 0.1
+ pbswgs = 0.79644 xrcrg1 = 12 xrcrg2 = 1
+ rbpb = 50 rbpd = 50 rbps = 50
+ rbdb = 50 rbsb = 50 gbmin = 1E-12
+ tnom = 30 ute = -0.9873002875 lute = -3.594247369143748E-7
+ kt1 = -0.25364 kt1l = 0 kt2 = -0.0391336648
+ lkt2 = 1.872936771156001E-8 ua1 = 2.119351845E-9 lua1 = 2.23825371687225E-15
+ ub1 = -1.1357150875E-18 lub1 = -5.198892232854376E-24 uc1 = -3.884688124999992E-12
+ luc1 = -6.098436109940627E-17 at = 6.113945334500001E5 lat = -1.106564669270528
+ prt = 0 njs = 1.2928 xtis = 2
+ tpb = 1.2287E-3 tpbsw = 0 tpbswg = 0
+ tcj = 7.92E-4 tcjsw = 1E-5 tcjswg = 0
+ tvoff = 0 tvfbsdoff = 0 saref = 3E-6
+ sbref = 3E-6 wlod = 0 ku0 = -2.7E-8
+ kvsat = 0.2 kvth0 = 7.9E-9 tku0 = 0
+ llodku0 = 0 wlodku0 = 1 llodvth = 0
+ wlodvth = 1 lku0 = 0 wku0 = 0
+ pku0 = 0 lkvth0 = 0 wkvth0 = 3E-7
+ pkvth0 = 0 stk2 = 0 lodk2 = 1
+ steta0 = 0 lodeta0 = 1

.model nlowvt_model.4 nmos
+ level = 54 lmin = 1E-6 lmax = 2E-6 wmin = 7E-6
+ wmax = 1.01E-3 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 4.148E-9
+ toxm = 4.148E-9 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 9.999999999999999E22 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {2.6E-8+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {1.2025E-8-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = -1.33E-8 dwb = -1.08E-8 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = 0.428149984201 lvth0 = 6.407049093034035E-9
+ vfb = 0 k1 = 0.4290139105 lk1 = 2.719084047525043E-9
+ k2 = -0.014261084845 lk2 = -7.993142885522248E-9 k3 = 1.65
+ k3b = 1.6 w0 = 1E-7 lpe0 = 2.3802E-7
+ lpeb = -4.9152E-8 vbm = -3 dvtp0 = 0
+ dvtp1 = 0 dvt0 = 0.07665 dvt1 = 0.1252
+ dvt2 = -0.05637 dvt0w = 0 dvt1w = 5.3E6
+ dvt2w = -0.032 vfbsdoff = 0 u0 = 0.038241159505
+ lu0 = -8.13391815890475E-9 ua = -9.501342297875E-10 lua = -5.427286937788895E-16
+ ub = 2.6177065205E-18 lub = 1.49665328318025E-25 uc = 5.966524835E-11
+ luc = 2.624012527281751E-17 ud = 0 up = 0
+ lp = 1 eu = 1.67 vsat = 1.918426775000001E4
+ lvsat = 0.051980787589387 a0 = 2.19057441012 la0 = -4.334906492266136E-7
+ ags = 0.81705744985 lags = 1.302146209218893E-6 b0 = 0
+ b1 = 0 keta = -0.1449161895 lketa = -7.827490885747496E-8
+ a1 = 0 a2 = 0.38689047 rdsw = 103.65
+ rdswmin = 0 rdw = 0 rdwmin = 0
+ rsw = 0 rswmin = 0 prwb = 0
+ prwg = 0 wr = 1 voff = -0.1170681977345
+ lvoff = 2.315097581485278E-9 voffl = 0 minv = 0
+ nfactor = 0.933140522895 lnfactor = 8.177035889556245E-7 eta0 = 5.91212287E-4
+ leta0 = -1.8023091849765E-10 etab = -5.41594989E-4 letab = 8.218961851454998E-11
+ dsub = -0.051530160903 ldsub = 6.609625482802829E-7 cit = 1.487975E-5
+ lcit = -9.642142012499999E-12 cdsc = 3.8556E-37 cdscb = -1.1484E-4
+ cdscd = 4.7984E-6 pclm = 0.2292314045 lpclm = 1.716301278225003E-9
+ pdiblc1 = 0.39 pdiblc2 = 7.015305875E-3 lpdiblc2 = 3.31207578129375E-9
+ pdiblcb = 0 drout = 3.4946 pscbe1 = 4.5E8
+ pscbe2 = 1E-8 pvag = 0 delta = 0.01
+ fprout = 0 pdits = 1.4427E-15 pditsl = 0
+ pditsd = 0 lambda = 0 vtl = 0
+ lc = 0 xn = 0 alpha0 = 1.8659456156935E-4
+ lalpha0 = -1.201672640344571E-10 alpha1 = 0 beta0 = 21.1969507455
+ lbeta0 = 1.969118241792744E-7 aigbacc = 1 bigbacc = 0
+ cigbacc = 0 nigbacc = 1 aigbinv = 0.35
+ bigbinv = 0.03 cigbinv = 6E-3 eigbinv = 1.1
+ nigbinv = 3 aigc = 0.43 bigc = 0.054
+ cigc = 0.075 aigsd = 0.43 bigsd = 0.054
+ cigsd = 0.075 dlcig = 0 nigc = 1
+ poxedge = 1 pigcd = 1 ntox = 1
+ toxref = 4.148E-9 agidl = 0 bgidl = 2.3E9
+ cgidl = 0.5 egidl = 0.8 noia = 9E41
+ noib = 1E27 noic = 8E11 em = 4.1E7
+ af = 1 ef = 1.2 kf = 0
+ lintnoi = -3E-7 tnoia = 2.5E7 tnoib = 9.9E6
+ ntnoi = 1 rnoia = 0.912 rnoib = 0.26
+ xpart = 0 cgso = {2.392894381E-10/sw_func_tox_lv_ratio} cgdo = {2.392894381E-10/sw_func_tox_lv_ratio}
+ cgbo = {1E-14/sw_func_tox_lv_ratio} ckappas = 0.6 cf = 1E-14
+ clc = 1E-7 cle = 0.6 dlc = 1.21071E-8
+ dwc = 2.6E-8 vfbcv = -1 noff = 3.8661
+ voffcv = -0.16994 acde = 0.38008 moin = 23.81
+ cgsl = {2.310725E-11/sw_func_tox_lv_ratio} cgdl = {2.310725E-11/sw_func_tox_lv_ratio} ijthsrev = 0.1
+ ijthsfwd = 0.1 xjbvs = 1 bvs = 11.9
+ jss = 2.75E-3 jsws = 6E-10 cjs = {1.210E-03*sw_func_nsd_pw_cj}
+ mjs = 0.42197 mjsws = 1E-3 cjsws = {3.230311424E-11*sw_func_nsd_pw_cj}
+ cjswgs = {1.795291232E-10*sw_func_nsd_pw_cj} mjswgs = 0.8 pbs = 0.7477
+ pbsws = 0.1 pbswgs = 0.79644 xrcrg1 = 12
+ xrcrg2 = 1 rbpb = 50 rbpd = 50
+ rbps = 50 rbdb = 50 rbsb = 50
+ gbmin = 1E-12 tnom = 30 ute = -1.32437605
+ lute = 3.066201159975E-7 kt1 = -0.250682631 lkt1 = -5.823853775549936E-9
+ kt1l = 0 kt2 = -0.04595043715 lkt2 = 3.219896903654249E-8
+ ua1 = 3.27396128E-9 lua1 = -4.319679621599968E-17 ub1 = -3.90831275E-18
+ lub1 = 2.796221183624992E-25 uc1 = 1.12738982E-11 luc1 = -9.093696974829E-17
+ at = 3.09962602E4 lat = 0.04027329875781 prt = 0
+ njs = 1.2928 xtis = 2 tpb = 1.2287E-3
+ tpbsw = 0 tpbswg = 0 tcj = 7.92E-4
+ tcjsw = 1E-5 tcjswg = 0 tvoff = 0
+ tvfbsdoff = 0 saref = 3E-6 sbref = 3E-6
+ wlod = 0 ku0 = -2.7E-8 kvsat = 0.2
+ kvth0 = 7.9E-9 tku0 = 0 llodku0 = 0
+ wlodku0 = 1 llodvth = 0 wlodvth = 1
+ lku0 = 0 wku0 = 0 pku0 = 0
+ lkvth0 = 0 wkvth0 = 3E-7 pkvth0 = 0
+ stk2 = 0 lodk2 = 1 steta0 = 0
+ lodeta0 = 1

.model nlowvt_model.5 nmos
+ level = 54 lmin = 5E-7 lmax = 1E-6 wmin = 7E-6
+ wmax = 1.01E-3 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 4.148E-9
+ toxm = 4.148E-9 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 9.999999999999999E22 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {2.6E-8+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {1.2025E-8-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = -1.33E-8 dwb = -1.08E-8 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = 0.441541299508 lvth0 = -6.662205080832581E-9
+ vfb = 0 k1 = 0.43379899 lk1 = -1.950914290499991E-9
+ k2 = -0.0171879335782 lk2 = -5.136684864355709E-9 k3 = 1.65
+ k3b = 1.6 w0 = 1E-7 lpe0 = 2.3802E-7
+ lpeb = -4.9152E-8 vbm = -3 dvtp0 = 0
+ dvtp1 = 0 dvt0 = 0.07665 dvt1 = 0.1252
+ dvt2 = -0.05637 dvt0w = 0 dvt1w = 5.3E6
+ dvt2w = -0.032 vfbsdoff = 0 u0 = 0.03407221921
+ lu0 = -4.065240877999501E-9 ua = -1.22160263213E-9 lua = -2.777891065127263E-16
+ ub = 2.751298556E-18 lub = 1.928618127179981E-26 uc = 1.074233594E-10
+ luc = -2.036940320643E-17 ud = 0 up = 0
+ lp = 1 eu = 1.67 vsat = 1.761046784000001E4
+ lvsat = 0.053516737611552 a0 = 2.02064512266 la0 = -2.676481611300271E-7
+ ags = 2.933555804800001 lags = -7.634503602945602E-7 b0 = 0
+ b1 = 0 keta = -0.43050084731601 lketa = 2.004414379380599E-7
+ a1 = 0 a2 = 0.38689047 rdsw = 103.65
+ rdswmin = 0 rdw = 0 rdwmin = 0
+ rsw = 0 rswmin = 0 prwb = 0
+ prwg = 0 wr = 1 voff = -0.114969616541
+ lvoff = 2.669872656889485E-10 voffl = 0 minv = 0
+ nfactor = 1.34690391681 lnfactor = 4.138912046642804E-7 eta0 = 7.840064259999999E-4
+ leta0 = -3.683883584546999E-10 etab = -8.332985404580999E-4 letab = 3.668776995600826E-10
+ dsub = 0.269443375494 ldsub = 3.477084254336306E-7 cit = 5E-6
+ cdsc = 3.8556E-37 cdscb = -1.1484E-4 cdscd = 4.7984E-6
+ pclm = -0.041272438 lpclm = 2.657145263660999E-7 pdiblc1 = 0.39
+ pdiblc2 = 0.0103033391 lpdiblc2 = 1.03119755355E-10 pdiblcb = 0
+ drout = 3.4946 pscbe1 = 4.5E8 pscbe2 = 1E-8
+ pvag = 0 delta = 0.01 fprout = 0
+ pdits = 1.4427E-15 pditsl = 0 pditsd = 0
+ lambda = 0 vtl = 0 lc = 0
+ xn = 0 alpha0 = -2.81603368637E-5 lalpha0 = 8.9422779091278E-11
+ alpha1 = 0 beta0 = 18.5608612212 lbeta0 = 2.76960339541986E-6
+ aigbacc = 1 bigbacc = 0 cigbacc = 0
+ nigbacc = 1 aigbinv = 0.35 bigbinv = 0.03
+ cigbinv = 6E-3 eigbinv = 1.1 nigbinv = 3
+ aigc = 0.43 bigc = 0.054 cigc = 0.075
+ aigsd = 0.43 bigsd = 0.054 cigsd = 0.075
+ dlcig = 0 nigc = 1 poxedge = 1
+ pigcd = 1 ntox = 1 toxref = 4.148E-9
+ agidl = 0 bgidl = 2.3E9 cgidl = 0.5
+ egidl = 0.8 noia = 9E41 noib = 1E27
+ noic = 8E11 em = 4.1E7 af = 1
+ ef = 1.2 kf = 0 lintnoi = -3E-7
+ tnoia = 2.5E7 tnoib = 9.9E6 ntnoi = 1
+ rnoia = 0.912 rnoib = 0.26 xpart = 0
+ cgso = {2.392894381E-10/sw_func_tox_lv_ratio} cgdo = {2.392894381E-10/sw_func_tox_lv_ratio} cgbo = {1E-14/sw_func_tox_lv_ratio}
+ ckappas = 0.6 cf = 1E-14 clc = 1E-7
+ cle = 0.6 dlc = 1.21071E-8 dwc = 2.6E-8
+ vfbcv = -1 noff = 3.8661 voffcv = -0.16994
+ acde = 0.38008 moin = 23.81 cgsl = {2.310725E-11/sw_func_tox_lv_ratio}
+ cgdl = {2.310725E-11/sw_func_tox_lv_ratio} ijthsrev = 0.1 ijthsfwd = 0.1
+ xjbvs = 1 bvs = 11.9 jss = 2.75E-3
+ jsws = 6E-10 cjs = {1.210E-03*sw_func_nsd_pw_cj} mjs = 0.42197
+ mjsws = 1E-3 cjsws = {3.230311424E-11*sw_func_nsd_pw_cj} cjswgs = {1.795291232E-10*sw_func_nsd_pw_cj}
+ mjswgs = 0.8 pbs = 0.7477 pbsws = 0.1
+ pbswgs = 0.79644 xrcrg1 = 12 xrcrg2 = 1
+ rbpb = 50 rbpd = 50 rbps = 50
+ rbdb = 50 rbsb = 50 gbmin = 1E-12
+ tnom = 30 ute = -1.00505974 lute = -5.016636747000065E-9
+ kt1 = -0.250681587 lkt1 = -5.824872667349997E-9 kt1l = 0
+ kt2 = -1.336252900000005E-3 lkt2 = -1.1342244082245E-8 ua1 = 4.02986714E-9
+ lua1 = -7.80923120283E-16 ub1 = -4.68630977E-18 lub1 = 1.0389083100315E-24
+ uc1 = -1.6803610036E-10 luc1 = 8.406062334634199E-17 at = 7.23638533E4
+ lat = -9.940372813499998E-5 prt = 0 njs = 1.2928
+ xtis = 2 tpb = 1.2287E-3 tpbsw = 0
+ tpbswg = 0 tcj = 7.92E-4 tcjsw = 1E-5
+ tcjswg = 0 tvoff = 0 tvfbsdoff = 0
+ saref = 2.74E-6 sbref = 2.74E-6 wlod = 0
+ ku0 = -2.7E-8 kvsat = 0.2 kvth0 = 7.9E-9
+ tku0 = 0 llodku0 = 0 wlodku0 = 1
+ llodvth = 0 wlodvth = 1 lku0 = 0
+ wku0 = 0 pku0 = 0 lkvth0 = 0
+ wkvth0 = 3E-7 pkvth0 = 0 stk2 = 0
+ lodk2 = 1 steta0 = 0 lodeta0 = 1

.model nlowvt_model.6 nmos
+ level = 54 lmin = 2.5E-7 lmax = 5E-7 wmin = 7E-6
+ wmax = 1.01E-3 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 4.148E-9
+ toxm = 4.148E-9 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 9.999999999999999E22 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {2.6E-8+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {1.2025E-8-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = -1.33E-8 dwb = -1.08E-8 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = 0.49556593788 lvth0 = -3.2375231713986E-8
+ vfb = 0 k1 = 0.29394924 lk1 = 6.461057422199998E-8
+ k2 = 0.0141190465532 lk2 = -2.003724205789553E-8 k3 = 1.65
+ k3b = 1.6 w0 = 1E-7 lpe0 = 2.3802E-7
+ lpeb = -4.9152E-8 vbm = -3 dvtp0 = 0
+ dvtp1 = 0 dvt0 = 0.07665 dvt1 = 0.1252
+ dvt2 = -0.05637 dvt0w = 0 dvt1w = 5.3E6
+ dvt2w = -0.032 vfbsdoff = 0 u0 = 0.027855798968
+ lu0 = -1.1065356638196E-9 ua = -1.68563919102E-9 lua = -5.693090630903107E-17
+ ub = 2.816927564E-18 lub = -1.194994508580004E-26 uc = 7.395486362740001E-11
+ luc = -4.440072643461033E-18 ud = 0 up = 0
+ lp = 1 eu = 1.67 vsat = 9.862158909799998E4
+ lvsat = 0.014959494448807 a0 = 1.31830138 la0 = 6.663234318900001E-8
+ ags = 2.5311021 lags = -5.719025194949999E-7 b0 = 0
+ b1 = 0 keta = -0.01362724653614 lketa = 2.030447646880833E-9
+ a1 = 0 a2 = 0.38689047 rdsw = 103.65
+ rdswmin = 0 rdw = 0 rdwmin = 0
+ rsw = 0 rswmin = 0 prwb = 0
+ prwg = 0 wr = 1 voff = -0.11864223996
+ lvoff = 2.014972381962E-9 voffl = 0 minv = 0
+ nfactor = 1.9844991982 lnfactor = 1.1042773048671E-7 eta0 = -5.197693882780001E-3
+ leta0 = 2.478601903509141E-9 etab = 0.024555479522316 letab = -1.171691121941734E-8
+ dsub = 1.659631036916 ldsub = -3.139513920201702E-7 cit = 5E-6
+ cdsc = 3.8556E-37 cdscb = -1.1484E-4 cdscd = 4.7984E-6
+ pclm = 0.640713106 lpclm = -5.887649330069999E-8 pdiblc1 = 0.39
+ pdiblc2 = 7.428100199999999E-3 lpdiblc2 = 1.47158970981E-9 pdiblcb = 0
+ drout = 3.4946 pscbe1 = 4.5E8 pscbe2 = 1E-8
+ pvag = 0 delta = 0.01 fprout = 0
+ pdits = 1.4427E-15 pditsl = 0 pditsd = 0
+ lambda = 0 vtl = 0 lc = 0
+ xn = 0 alpha0 = -2.283466401976E-3 lalpha0 = 1.162835700781477E-9
+ alpha1 = 0 beta0 = 18.1542346952 lbeta0 = 2.96313729046956E-6
+ aigbacc = 1 bigbacc = 0 cigbacc = 0
+ nigbacc = 1 aigbinv = 0.35 bigbinv = 0.03
+ cigbinv = 6E-3 eigbinv = 1.1 nigbinv = 3
+ aigc = 0.43 bigc = 0.054 cigc = 0.075
+ aigsd = 0.43 bigsd = 0.054 cigsd = 0.075
+ dlcig = 0 nigc = 1 poxedge = 1
+ pigcd = 1 ntox = 1 toxref = 4.148E-9
+ agidl = 0 bgidl = 2.3E9 cgidl = 0.5
+ egidl = 0.8 noia = 9E41 noib = 1E27
+ noic = 8E11 em = 4.1E7 af = 1
+ ef = 1.2 kf = 0 lintnoi = -3E-7
+ tnoia = 2.5E7 tnoib = 9.9E6 ntnoi = 1
+ rnoia = 0.912 rnoib = 0.26 xpart = 0
+ cgso = {2.392894381E-10/sw_func_tox_lv_ratio} cgdo = {2.392894381E-10/sw_func_tox_lv_ratio} cgbo = {1E-14/sw_func_tox_lv_ratio}
+ ckappas = 0.6 cf = 1E-14 clc = 1E-7
+ cle = 0.6 dlc = 1.21071E-8 dwc = 2.6E-8
+ vfbcv = -1 noff = 3.8661 voffcv = -0.16994
+ acde = 0.38008 moin = 23.81 cgsl = {2.310725E-11/sw_func_tox_lv_ratio}
+ cgdl = {2.310725E-11/sw_func_tox_lv_ratio} ijthsrev = 0.1 ijthsfwd = 0.1
+ xjbvs = 1 bvs = 11.9 jss = 2.75E-3
+ jsws = 6E-10 cjs = {1.210E-03*sw_func_nsd_pw_cj} mjs = 0.42197
+ mjsws = 1E-3 cjsws = {3.230311424E-11*sw_func_nsd_pw_cj} cjswgs = {1.795291232E-10*sw_func_nsd_pw_cj}
+ mjswgs = 0.8 pbs = 0.7477 pbsws = 0.1
+ pbswgs = 0.79644 xrcrg1 = 12 xrcrg2 = 1
+ rbpb = 50 rbpd = 50 rbps = 50
+ rbdb = 50 rbsb = 50 gbmin = 1E-12
+ tnom = 30 ute = -0.4267743 lute = -2.80251591915E-7
+ kt1 = -0.253945266 lkt1 = -4.271524647299997E-9 kt1l = 0
+ kt2 = -0.0283510874 lkt2 = 1.515466398029999E-9 ua1 = 4.105298706E-9
+ lua1 = -8.168247741206999E-16 ub1 = -4.131849346E-18 lub1 = 7.750128712286998E-25
+ uc1 = 4.935840992E-11 luc1 = -1.9408293821424E-17 at = 8.74644682E4
+ lat = -7.286541389789999E-3 prt = 0 njs = 1.2928
+ xtis = 2 tpb = 1.2287E-3 tpbsw = 0
+ tpbswg = 0 tcj = 7.92E-4 tcjsw = 1E-5
+ tcjswg = 0 tvoff = 0 tvfbsdoff = 0
+ saref = 1.74E-6 sbref = 1.74E-6 wlod = 0
+ ku0 = -2.7E-8 kvsat = 0.2 kvth0 = 7.9E-9
+ tku0 = 0 llodku0 = 0 wlodku0 = 1
+ llodvth = 0 wlodvth = 1 lku0 = 0
+ wku0 = 0 pku0 = 0 lkvth0 = 0
+ wkvth0 = 3E-7 pkvth0 = 0 stk2 = 0
+ lodk2 = 1 steta0 = 0 lodeta0 = 1

.model nlowvt_model.7 nmos
+ level = 54 lmin = 1.8E-7 lmax = 2.5E-7 wmin = 7E-6
+ wmax = 1.01E-3 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 4.148E-9
+ toxm = 4.148E-9 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 9.999999999999999E22 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {2.6E-8+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {1.2025E-8-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = -1.33E-8 dwb = -1.08E-8 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = 0.608598192142857 lvth0 = -5.791486956467857E-8
+ vfb = 0 k1 = 0.315631585714286 lk1 = 5.971144820785717E-8
+ k2 = -4.315366052857122E-3 lk2 = -1.587198652955693E-8 k3 = 1.65
+ k3b = 1.6 w0 = 1E-7 lpe0 = 2.3802E-7
+ lpeb = -4.9152E-8 vbm = -3 dvtp0 = 0
+ dvtp1 = 0 dvt0 = 0.07665 dvt1 = 0.1252
+ dvt2 = -0.05637 dvt0w = 0 dvt1w = 5.3E6
+ dvt2w = -0.032 vfbsdoff = 0 u0 = 0.03935215995
+ lu0 = -3.704138427702499E-9 ua = -9.341333047142863E-10 lua = -2.26733661319807E-16
+ ub = 2.603968464285714E-18 lub = 3.616816349464292E-26 uc = 8.319096704499999E-11
+ luc = -6.526970210667748E-18 ud = 0 up = 0
+ lp = 1 eu = 1.67 vsat = 1.521236440071429E5
+ lvsat = 2.87070514208607E-3 a0 = 5.207179142857143 la0 = -8.120595873285714E-7
+ ags = -2.681894428571429 lags = 6.059740461357142E-7 b0 = 0
+ b1 = 0 keta = 0.246367573079143 lketa = -5.671538184519232E-8
+ a1 = 0 a2 = 0.38689047 rdsw = 103.65
+ rdswmin = 0 rdw = 0 rdwmin = 0
+ rsw = 0 rswmin = 0 prwb = 0
+ prwg = 0 wr = 1 voff = -0.163941736239286
+ lvoff = 1.22503935662666E-8 voffl = 0 minv = 0
+ nfactor = 1.251539365928572 lnfactor = 2.760400045884392E-7 eta0 = -0.153900091517214
+ leta0 = 3.607790864900957E-8 etab = -0.055089748665714 letab = 6.278928089668142E-9
+ dsub = 0.154872654907143 ldsub = 2.604876439473105E-8 cit = 5E-6
+ cdsc = 3.8556E-37 cdscb = -1.1484E-4 cdscd = 4.7984E-6
+ pclm = 0.896579564285714 lpclm = -1.166895195503571E-7 pdiblc1 = -0.968992857142857
+ lpdiblc1 = 3.070644360714285E-7 pdiblc2 = 0.014460090714286 lpdiblc2 = -1.172885468928574E-10
+ pdiblcb = 0 drout = 3.4946 pscbe1 = 4.5E8
+ pscbe2 = 1E-8 pvag = 0 delta = 0.01
+ fprout = 0 pdits = 1.4427E-15 pditsl = 0
+ pditsd = 0 lambda = 0 vtl = 0
+ lc = 0 xn = 0 alpha0 = 7.807445427571428E-3
+ lalpha0 = -1.117205827104764E-9 alpha1 = 0 beta0 = 36.324204075714285
+ lbeta0 = -1.142367291057642E-6 aigbacc = 1 bigbacc = 0
+ cigbacc = 0 nigbacc = 1 aigbinv = 0.35
+ bigbinv = 0.03 cigbinv = 6E-3 eigbinv = 1.1
+ nigbinv = 3 aigc = 0.43 bigc = 0.054
+ cigc = 0.075 aigsd = 0.43 bigsd = 0.054
+ cigsd = 0.075 dlcig = 0 nigc = 1
+ poxedge = 1 pigcd = 1 ntox = 1
+ toxref = 4.148E-9 agidl = 0 bgidl = 2.3E9
+ cgidl = 0.5 egidl = 0.8 noia = 9E41
+ noib = 1E27 noic = 8E11 em = 4.1E7
+ af = 1 ef = 1.2 kf = 0
+ lintnoi = -3E-7 tnoia = 2.5E7 tnoib = 9.9E6
+ ntnoi = 1 rnoia = 0.912 rnoib = 0.26
+ xpart = 0 cgso = {2.392894381E-10/sw_func_tox_lv_ratio} cgdo = {2.392894381E-10/sw_func_tox_lv_ratio}
+ cgbo = {1E-14/sw_func_tox_lv_ratio} ckappas = 0.6 cf = 1E-14
+ clc = 1E-7 cle = 0.6 dlc = 1.21071E-8
+ dwc = 2.6E-8 vfbcv = -1 noff = 3.8661
+ voffcv = -0.16994 acde = 0.38008 moin = 23.81
+ cgsl = {2.310725E-11/sw_func_tox_lv_ratio} cgdl = {2.310725E-11/sw_func_tox_lv_ratio} ijthsrev = 0.1
+ ijthsfwd = 0.1 xjbvs = 1 bvs = 11.9
+ jss = 2.75E-3 jsws = 6E-10 cjs = {1.210E-03*sw_func_nsd_pw_cj}
+ mjs = 0.42197 mjsws = 1E-3 cjsws = {3.230311424E-11*sw_func_nsd_pw_cj}
+ cjswgs = {1.795291232E-10*sw_func_nsd_pw_cj} mjswgs = 0.8 pbs = 0.7477
+ pbsws = 0.1 pbswgs = 0.79644 xrcrg1 = 12
+ xrcrg2 = 1 rbpb = 50 rbpd = 50
+ rbps = 50 rbdb = 50 rbsb = 50
+ gbmin = 1E-12 tnom = 30 ute = -1.139543428571429
+ lute = -1.192014073142856E-7 kt1 = -0.182176214285714 lkt1 = -2.048774188214286E-8
+ kt1l = 0 kt2 = -0.035109168571429 lkt2 = 3.042454838714286E-9
+ ua1 = 1.54170728E-9 lua1 = -2.37581291416E-16 ub1 = -1.9959031E-18
+ lub1 = 2.92395816945E-25 uc1 = -1.221356132142857E-10 luc1 = 1.934078070576786E-17
+ at = 136.68785714285332 lat = 0.012445170578679 prt = 0
+ njs = 1.2928 xtis = 2 tpb = 1.2287E-3
+ tpbsw = 0 tpbswg = 0 tcj = 7.92E-4
+ tcjsw = 1E-5 tcjswg = 0 tvoff = 0
+ tvfbsdoff = 0 saref = 1.25E-6 sbref = 1.24E-6
+ wlod = 0 ku0 = -2.7E-8 kvsat = 0.2
+ kvth0 = 7.9E-9 tku0 = 0 llodku0 = 0
+ wlodku0 = 1 llodvth = 0 wlodvth = 1
+ lku0 = 0 wku0 = 0 pku0 = 0
+ lkvth0 = 0 wkvth0 = 3E-7 pkvth0 = 0
+ stk2 = 0 lodk2 = 1 steta0 = 0
+ lodeta0 = 1

.model nlowvt_model.8 nmos
+ level = 54 lmin = 1.5E-7 lmax = 1.8E-7 wmin = 7E-6
+ wmax = 1.01E-3 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 4.148E-9
+ toxm = 4.148E-9 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 9.999999999999999E22 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {2.6E-8+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {1.2025E-8-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = -1.33E-8 dwb = -1.08E-8 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = 0.249959346666667 lvth0 = -1.985141612666671E-9
+ vfb = 0 k1 = 1.011211866666667 lk1 = -4.876429660666666E-8
+ k2 = -0.21737859252 lk2 = 1.7355223637994E-8 k3 = 1.65
+ k3b = 1.6 w0 = 1E-7 lpe0 = 2.3802E-7
+ lpeb = -4.9152E-8 vbm = -3 dvtp0 = 0
+ dvtp1 = 0 dvt0 = 0.07665 dvt1 = 0.1252
+ dvt2 = -0.05637 dvt0w = 0 dvt1w = 5.3E6
+ dvt2w = -0.032 vfbsdoff = 0 u0 = 0.01421071555
+ lu0 = 2.166698264775001E-10 ua = -3.496851672833332E-9 lua = 1.729222681883582E-16
+ ub = 4.57941585E-18 lub = -2.719028563075E-25 uc = 1.863698448333334E-10
+ luc = -2.261771620175834E-17 ud = 0 up = 0
+ lp = 1 eu = 1.67 vsat = 1.819855189500001E5
+ lvsat = -1.786254255252507E-3 a0 = 0 ags = 1.005218833333333
+ lags = 3.096873294166675E-8 b0 = 0 b1 = 0
+ keta = 0.1569286063 lketa = -4.276737497598501E-8 a1 = 0
+ a2 = 0.38689047 rdsw = 103.65 rdswmin = 0
+ rdw = 0 rdwmin = 0 rsw = 0
+ rswmin = 0 prwb = 0 prwg = 0
+ wr = 1 voff = -0.11934831869 lvoff = 5.296050099455504E-9
+ voffl = 0 minv = 0 nfactor = 0.723459400166666
+ lnfactor = 3.583940752490084E-7 eta0 = 0.067637351756667 leta0 = 1.529144370447834E-9
+ etab = -0.077077273825 letab = 9.70788263825875E-9 dsub = 0.58180516425
+ ldsub = -4.053136043728748E-8 cit = 5E-6 cdsc = 3.8556E-37
+ cdscb = -1.1484E-4 cdscd = 4.7984E-6 pclm = 0.086824416666667
+ lpclm = 9.59179572083335E-9 pdiblc1 = 3.583688213883334 lpdiblc1 = -4.029261769551058E-7
+ pdiblc2 = 0.064735802833333 lpdiblc2 = -7.957785851858334E-9 pdiblcb = 0
+ drout = 3.4946 pscbe1 = 4.5E8 pscbe2 = 1E-8
+ pvag = 0 delta = 0.01 fprout = 0
+ pdits = 1.4427E-15 pditsl = 0 pditsd = 0
+ lambda = 0 vtl = 0 lc = 0
+ xn = 0 alpha0 = 1.687407635666667E-3 lalpha0 = -1.627859334572167E-10
+ alpha1 = 0 beta0 = 31.24083182666667 lbeta0 = -3.496153888186668E-7
+ aigbacc = 1 bigbacc = 0 cigbacc = 0
+ nigbacc = 1 aigbinv = 0.35 bigbinv = 0.03
+ cigbinv = 6E-3 eigbinv = 1.1 nigbinv = 3
+ aigc = 0.43 bigc = 0.054 cigc = 0.075
+ aigsd = 0.43 bigsd = 0.054 cigsd = 0.075
+ dlcig = 0 nigc = 1 poxedge = 1
+ pigcd = 1 ntox = 1 toxref = 4.148E-9
+ agidl = 0 bgidl = 2.3E9 cgidl = 0.5
+ egidl = 0.8 noia = 9E41 noib = 1E27
+ noic = 8E11 em = 4.1E7 af = 1
+ ef = 1.2 kf = 0 lintnoi = -3E-7
+ tnoia = 2.5E7 tnoib = 9.9E6 ntnoi = 1
+ rnoia = 0.912 rnoib = 0.26 xpart = 0
+ cgso = {2.392894381E-10/sw_func_tox_lv_ratio} cgdo = {2.392894381E-10/sw_func_tox_lv_ratio} cgbo = {1E-14/sw_func_tox_lv_ratio}
+ ckappas = 0.6 cf = 1E-14 clc = 1E-7
+ cle = 0.6 dlc = 1.21071E-8 dwc = 2.6E-8
+ vfbcv = -1 noff = 3.8661 voffcv = -0.16994
+ acde = 0.38008 moin = 23.81 cgsl = {2.310725E-11/sw_func_tox_lv_ratio}
+ cgdl = {2.310725E-11/sw_func_tox_lv_ratio} ijthsrev = 0.1 ijthsfwd = 0.1
+ xjbvs = 1 bvs = 11.9 jss = 2.75E-3
+ jsws = 6E-10 cjs = {1.210E-03*sw_func_nsd_pw_cj} mjs = 0.42197
+ mjsws = 1E-3 cjsws = {3.230311424E-11*sw_func_nsd_pw_cj} cjswgs = {1.795291232E-10*sw_func_nsd_pw_cj}
+ mjswgs = 0.8 pbs = 0.7477 pbsws = 0.1
+ pbswgs = 0.79644 xrcrg1 = 12 xrcrg2 = 1
+ rbpb = 50 rbpd = 50 rbps = 50
+ rbdb = 50 rbsb = 50 gbmin = 1E-12
+ tnom = 30 ute = -2.841387833333333 lute = 1.462012276083332E-7
+ kt1 = -0.295119316666667 lkt1 = -2.874265065833337E-9 kt1l = 0
+ kt2 = 0.02122778 lkt2 = -5.743292291000001E-9 ua1 = -2.42902207E-9
+ lua1 = 3.816539507165E-16 ub1 = 2.4443796E-18 lub1 = -4.0006627012E-25
+ uc1 = 5.2148775E-12 luc1 = -5.195283211249999E-19 at = 6.394335E4
+ lat = 2.4945216175E-3 prt = 0 njs = 1.2928
+ xtis = 2 tpb = 1.2287E-3 tpbsw = 0
+ tpbswg = 0 tcj = 7.92E-4 tcjsw = 1E-5
+ tcjswg = 0 tvoff = 0 tvfbsdoff = 0
+ saref = 1.1E-6 sbref = 1.1E-6 wlod = 0
+ ku0 = -2.7E-8 kvsat = 0.2 kvth0 = 7.9E-9
+ tku0 = 0 llodku0 = 0 wlodku0 = 1
+ llodvth = 0 wlodvth = 1 lku0 = 0
+ wku0 = 0 pku0 = 0 lkvth0 = 0
+ wkvth0 = 3E-7 pkvth0 = 0 stk2 = 0
+ lodk2 = 1 steta0 = 0 lodeta0 = 1

.model nlowvt_model.9 nmos
+ level = 54 lmin = 8E-6 lmax = 2.02E-5 wmin = 5E-6
+ wmax = 7E-6 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 4.148E-9
+ toxm = 4.148E-9 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 9.999999999999999E22 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {2.6E-8+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {1.2025E-8-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = -1.33E-8 dwb = -1.08E-8 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = 0.3916346148 wvth0 = 1.825474803696003E-7
+ vfb = 0 k1 = 0.64981268 wk1 = -1.23453926064E-6
+ k2 = -0.094489771866 wk2 = 4.252715989249682E-7 k3 = 1.65
+ k3b = 1.6 w0 = 1E-7 lpe0 = 2.3802E-7
+ lpeb = -4.9152E-8 vbm = -3 dvtp0 = 0
+ dvtp1 = 0 dvt0 = 0.07665 dvt1 = 0.1252
+ dvt2 = -0.05637 dvt0w = 0 dvt1w = 5.3E6
+ dvt2w = -0.032 vfbsdoff = 0 u0 = 0.03097422792
+ wu0 = 7.046259171840022E-9 ua = -1.3902455543E-9 wua = 6.161858416764019E-16
+ ub = 2.711605659999999E-18 wub = -2.507926456799964E-25 uc = 6.9437014E-11
+ wuc = 4.967722727999962E-18 ud = 0 up = 0
+ lp = 1 eu = 1.67 vsat = -4.125794000000012E4
+ wvsat = 1.406260887120001 a0 = 2.0466021424 wa0 = -6.027893201952018E-7
+ ags = 0.4928656944 wags = 2.704641401088007E-7 b0 = 0
+ b1 = 0 keta = 0 a1 = 0
+ a2 = 0.38689047 rdsw = 103.65 rdswmin = 0
+ rdw = 0 rdwmin = 0 rsw = 0
+ rswmin = 0 prwb = 0 prwg = 0
+ wr = 1 voff = -0.10742454972 wvoff = -5.679740066543997E-8
+ voffl = 0 minv = 0 nfactor = 1.30077583784
+ wnfactor = -1.381734432112321E-6 eta0 = 0.08 etab = -0.07
+ dsub = 0.56 cit = 1E-5 cdsc = 3.8556E-37
+ cdscb = -1.1484E-4 cdscd = 4.7984E-6 pclm = 0.525464596
+ wpclm = -2.261328013008001E-6 pdiblc1 = 0.39 pdiblc2 = 3.709717999999989E-4
+ wpdiblc2 = 3.075690753360001E-8 pdiblcb = 0 drout = 3.4946
+ pscbe1 = 4.5E8 pscbe2 = 1E-8 pvag = 0
+ delta = 0.01 fprout = 0 pdits = 1.4427E-15
+ pditsl = 0 pditsd = 0 lambda = 0
+ vtl = 0 lc = 0 xn = 0
+ alpha0 = 2.094204810660001E-4 walpha0 = -8.690198776105684E-10 alpha1 = 0
+ beta0 = 18.519724724 wbeta0 = -4.84096844635199E-6 aigbacc = 1
+ bigbacc = 0 cigbacc = 0 nigbacc = 1
+ aigbinv = 0.35 bigbinv = 0.03 cigbinv = 6E-3
+ eigbinv = 1.1 nigbinv = 3 aigc = 0.43
+ bigc = 0.054 cigc = 0.075 aigsd = 0.43
+ bigsd = 0.054 cigsd = 0.075 dlcig = 0
+ nigc = 1 poxedge = 1 pigcd = 1
+ ntox = 1 toxref = 4.148E-9 agidl = 0
+ bgidl = 2.3E9 cgidl = 0.5 egidl = 0.8
+ noia = 9E41 noib = 1E27 noic = 8E11
+ em = 4.1E7 af = 1 ef = 1.2
+ kf = 0 lintnoi = -3E-7 tnoia = 2.5E7
+ tnoib = 9.9E6 ntnoi = 1 rnoia = 0.912
+ rnoib = 0.26 xpart = 0 cgso = {2.392894381E-10/sw_func_tox_lv_ratio}
+ cgdo = {2.392894381E-10/sw_func_tox_lv_ratio} cgbo = {1E-14/sw_func_tox_lv_ratio} ckappas = 0.6
+ cf = 1E-14 clc = 1E-7 cle = 0.6
+ dlc = 1.21071E-8 dwc = 2.6E-8 vfbcv = -1
+ noff = 3.8661 voffcv = -0.16994 acde = 0.38008
+ moin = 23.81 cgsl = {2.310725E-11/sw_func_tox_lv_ratio} cgdl = {2.310725E-11/sw_func_tox_lv_ratio}
+ ijthsrev = 0.1 ijthsfwd = 0.1 xjbvs = 1
+ bvs = 11.9 jss = 2.75E-3 jsws = 6E-10
+ cjs = {1.210E-03*sw_func_nsd_pw_cj} mjs = 0.42197 mjsws = 1E-3
+ cjsws = {3.230311424E-11*sw_func_nsd_pw_cj} cjswgs = {1.795291232E-10*sw_func_nsd_pw_cj} mjswgs = 0.8
+ pbs = 0.7477 pbsws = 0.1 pbswgs = 0.79644
+ xrcrg1 = 12 xrcrg2 = 1 rbpb = 50
+ rbpd = 50 rbps = 50 rbdb = 50
+ rbsb = 50 gbmin = 1E-12 tnom = 30
+ ute = -0.7827992 wute = -2.0489707584E-6 kt1 = -0.25267514
+ wkt1 = -6.703847280000028E-9 kt1l = 0 kt2 = -0.033762442
+ wkt2 = -4.58955698399994E-9 ua1 = 2.081118E-9 wua1 = 4.177012535999996E-15
+ ub1 = -3.903747999999989E-19 wub1 = -1.426372428960001E-23 uc1 = -3.712999999999178E-14
+ wuc1 = -1.333034247600001E-16 at = 9.886528900000002E5 wat = -4.554920439720002
+ prt = 0 njs = 1.2928 xtis = 2
+ tpb = 1.2287E-3 tpbsw = 0 tpbswg = 0
+ tcj = 7.92E-4 tcjsw = 1E-5 tcjswg = 0
+ tvoff = 0 tvfbsdoff = 0 saref = 3E-6
+ sbref = 3E-6 wlod = 0 ku0 = -2.7E-8
+ kvsat = 0.2 kvth0 = 7.9E-9 tku0 = 0
+ llodku0 = 0 wlodku0 = 1 llodvth = 0
+ wlodvth = 1 lku0 = 0 wku0 = 0
+ pku0 = 0 lkvth0 = 0 wkvth0 = 3E-7
+ pkvth0 = 0 stk2 = 0 lodk2 = 1
+ steta0 = 0 lodeta0 = 1

.model nlowvt_model.10 nmos
+ level = 54 lmin = 4E-6 lmax = 8E-6 wmin = 5E-6
+ wmax = 7E-6 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 4.148E-9
+ toxm = 4.148E-9 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 9.999999999999999E22 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {2.6E-8+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {1.2025E-8-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = -1.33E-8 dwb = -1.08E-8 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = 0.3916346148 wvth0 = 1.825474803696003E-7
+ vfb = 0 k1 = 0.64981268 wk1 = -1.23453926064E-6
+ k2 = -0.094489771866 wk2 = 4.252715989249682E-7 k3 = 1.65
+ k3b = 1.6 w0 = 1E-7 lpe0 = 2.3802E-7
+ lpeb = -4.9152E-8 vbm = -3 dvtp0 = 0
+ dvtp1 = 0 dvt0 = 0.07665 dvt1 = 0.1252
+ dvt2 = -0.05637 dvt0w = 0 dvt1w = 5.3E6
+ dvt2w = -0.032 vfbsdoff = 0 u0 = 0.03097422792
+ wu0 = 7.046259171840022E-9 ua = -1.3902455543E-9 wua = 6.161858416764019E-16
+ ub = 2.711605659999999E-18 wub = -2.507926456799964E-25 uc = 6.9437014E-11
+ wuc = 4.967722727999962E-18 ud = 0 up = 0
+ lp = 1 eu = 1.67 vsat = -4.125794000000012E4
+ wvsat = 1.406260887120001 a0 = 2.0466021424 wa0 = -6.027893201952018E-7
+ ags = 0.4928656944 wags = 2.704641401088007E-7 b0 = 0
+ b1 = 0 keta = 0 a1 = 0
+ a2 = 0.38689047 rdsw = 103.65 rdswmin = 0
+ rdw = 0 rdwmin = 0 rsw = 0
+ rswmin = 0 prwb = 0 prwg = 0
+ wr = 1 voff = -0.10742454972 wvoff = -5.679740066543997E-8
+ voffl = 0 minv = 0 nfactor = 1.30077583784
+ wnfactor = -1.381734432112321E-6 eta0 = 0.08 etab = -0.07
+ dsub = 0.56 cit = 1E-5 cdsc = 3.8556E-37
+ cdscb = -1.1484E-4 cdscd = 4.7984E-6 pclm = 0.525464596
+ wpclm = -2.261328013008001E-6 pdiblc1 = 0.39 pdiblc2 = 3.709717999999989E-4
+ wpdiblc2 = 3.075690753360001E-8 pdiblcb = 0 drout = 3.4946
+ pscbe1 = 4.5E8 pscbe2 = 1E-8 pvag = 0
+ delta = 0.01 fprout = 0 pdits = 1.4427E-15
+ pditsl = 0 pditsd = 0 lambda = 0
+ vtl = 0 lc = 0 xn = 0
+ alpha0 = 2.094204810660001E-4 walpha0 = -8.690198776105684E-10 alpha1 = 0
+ beta0 = 18.519724724 wbeta0 = -4.84096844635199E-6 aigbacc = 1
+ bigbacc = 0 cigbacc = 0 nigbacc = 1
+ aigbinv = 0.35 bigbinv = 0.03 cigbinv = 6E-3
+ eigbinv = 1.1 nigbinv = 3 aigc = 0.43
+ bigc = 0.054 cigc = 0.075 aigsd = 0.43
+ bigsd = 0.054 cigsd = 0.075 dlcig = 0
+ nigc = 1 poxedge = 1 pigcd = 1
+ ntox = 1 toxref = 4.148E-9 agidl = 0
+ bgidl = 2.3E9 cgidl = 0.5 egidl = 0.8
+ noia = 9E41 noib = 1E27 noic = 8E11
+ em = 4.1E7 af = 1 ef = 1.2
+ kf = 0 lintnoi = -3E-7 tnoia = 2.5E7
+ tnoib = 9.9E6 ntnoi = 1 rnoia = 0.912
+ rnoib = 0.26 xpart = 0 cgso = {2.392894381E-10/sw_func_tox_lv_ratio}
+ cgdo = {2.392894381E-10/sw_func_tox_lv_ratio} cgbo = {1E-14/sw_func_tox_lv_ratio} ckappas = 0.6
+ cf = 1E-14 clc = 1E-7 cle = 0.6
+ dlc = 1.21071E-8 dwc = 2.6E-8 vfbcv = -1
+ noff = 3.8661 voffcv = -0.16994 acde = 0.38008
+ moin = 23.81 cgsl = {2.310725E-11/sw_func_tox_lv_ratio} cgdl = {2.310725E-11/sw_func_tox_lv_ratio}
+ ijthsrev = 0.1 ijthsfwd = 0.1 xjbvs = 1
+ bvs = 11.9 jss = 2.75E-3 jsws = 6E-10
+ cjs = {1.210E-03*sw_func_nsd_pw_cj} mjs = 0.42197 mjsws = 1E-3
+ cjsws = {3.230311424E-11*sw_func_nsd_pw_cj} cjswgs = {1.795291232E-10*sw_func_nsd_pw_cj} mjswgs = 0.8
+ pbs = 0.7477 pbsws = 0.1 pbswgs = 0.79644
+ xrcrg1 = 12 xrcrg2 = 1 rbpb = 50
+ rbpd = 50 rbps = 50 rbdb = 50
+ rbsb = 50 gbmin = 1E-12 tnom = 30
+ ute = -0.7827992 wute = -2.0489707584E-6 kt1 = -0.25267514
+ wkt1 = -6.703847280000028E-9 kt1l = 0 kt2 = -0.033762442
+ wkt2 = -4.58955698399994E-9 ua1 = 2.081118E-9 wua1 = 4.177012535999996E-15
+ ub1 = -3.903747999999989E-19 wub1 = -1.426372428960001E-23 uc1 = -3.712999999999178E-14
+ wuc1 = -1.333034247600001E-16 at = 9.886528900000002E5 wat = -4.554920439720002
+ prt = 0 njs = 1.2928 xtis = 2
+ tpb = 1.2287E-3 tpbsw = 0 tpbswg = 0
+ tcj = 7.92E-4 tcjsw = 1E-5 tcjswg = 0
+ tvoff = 0 tvfbsdoff = 0 saref = 3E-6
+ sbref = 3E-6 wlod = 0 ku0 = -2.7E-8
+ kvsat = 0.2 kvth0 = 7.9E-9 tku0 = 0
+ llodku0 = 0 wlodku0 = 1 llodvth = 0
+ wlodvth = 1 lku0 = 0 wku0 = 0
+ pku0 = 0 lkvth0 = 0 wkvth0 = 3E-7
+ pkvth0 = 0 stk2 = 0 lodk2 = 1
+ steta0 = 0 lodeta0 = 1

.model nlowvt_model.11 nmos
+ level = 54 lmin = 2E-6 lmax = 4E-6 wmin = 5E-6
+ wmax = 7E-6 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 4.148E-9
+ toxm = 4.148E-9 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 9.999999999999999E22 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {2.6E-8+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {1.2025E-8-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = -1.33E-8 dwb = -1.08E-8 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = 0.340996998785017 lvth0 = 2.013326293947703E-7
+ wvth0 = 4.418139563713496E-7 pvth0 = -1.030830545259155E-12 vfb = 0
+ k1 = 1.025228637008 lk1 = -1.492635074265958E-6 wk1 = -3.556407174409586E-6
+ pk1 = 9.231630731752184E-12 k2 = -0.228175449342856 lk2 = 5.315275693641072E-7
+ wk2 = 1.251319737676456E-6 pk2 = -3.28432609726898E-12 k3 = 1.65
+ k3b = 1.6 w0 = 1E-7 lpe0 = 2.3802E-7
+ lpeb = -4.9152E-8 vbm = -3 dvtp0 = 0
+ dvtp1 = 0 dvt0 = 0.07665 dvt1 = 0.1252
+ dvt2 = -0.05637 dvt0w = 0 dvt1w = 5.3E6
+ dvt2w = -0.032 vfbsdoff = 0 u0 = 0.024725202916783
+ lu0 = 2.484581096153869E-8 wu0 = 3.579975378478936E-8 pu0 = -1.143224569063559E-13
+ ua = -1.619441111917716E-9 lua = 9.112700773101556E-16 wua = 1.681729951539163E-15
+ pua = -4.236550103608845E-21 ub = 2.608797040778498E-18 lub = 4.087619295937291E-25
+ wub = 3.403734022889948E-25 pub = -2.35044664842231E-30 uc = 1.231031145377501E-10
+ luc = -2.133737324330673E-16 wuc = -3.870767534961874E-16 puc = 1.558749235243558E-21
+ ud = 0 up = 0 lp = 1
+ eu = 1.67 vsat = -1.193254422777502E5 lvsat = 0.31039248568122
+ wvsat = 2.742540705690509 pvsat = -5.312981744645411E-6 a0 = 1.996896517090061
+ la0 = 1.976270809510549E-7 wa0 = -3.353193750905698E-7 pa0 = -1.063447128238761E-12
+ ags = -0.66403401168606 lags = 4.59977538641287E-6 wags = 1.826760983036024E-6
+ pags = -6.187758432636494E-12 b0 = 0 b1 = 0
+ keta = 0.1053904745295 lketa = -4.190272572055656E-7 wketa = 5.344439968280344E-7
+ pketa = -2.124922609188423E-12 a1 = 0 a2 = 0.38689047
+ rdsw = 103.65 rdswmin = 0 rdw = 0
+ rdwmin = 0 rsw = 0 rswmin = 0
+ prwb = 0 prwg = 0 wr = 1
+ voff = -0.087942976394225 lvoff = -7.745776146461701E-8 wvoff = -1.901140905472171E-7
+ pvoff = 5.300604931354516E-13 voffl = 0 minv = 0
+ nfactor = 1.733084749283323 lnfactor = -1.718838616453079E-6 wnfactor = -6.067623744453739E-6
+ pnfactor = 1.863086161140386E-11 eta0 = 0.1585440125 leta0 = -3.122870664993751E-7
+ etab = -0.1386642625 letab = 2.730056744868751E-7 dsub = 1.17193790508545
+ ldsub = -2.433034513724496E-6 wdsub = -2.350110060789765E-6 pdsub = 9.343920096197066E-12
+ cit = -2.221250750000012E-6 lcit = 4.859108191946253E-11 wcit = 8.491325021100008E-11
+ pcit = -3.376108371764257E-16 cdsc = 3.8556E-37 cdscb = -1.1484E-4
+ cdscd = 4.7984E-6 pclm = 0.375371671114 lpclm = 5.967619647004922E-7
+ wpclm = -1.425102324930072E-6 ppclm = -3.324791524513441E-12 pdiblc1 = 0.39
+ pdiblc2 = -7.624875459610005E-3 lpdiblc2 = 3.179108891184638E-8 wpdiblc2 = 5.95832577152303E-8
+ ppdiblc2 = -1.146121270046529E-13 pdiblcb = 0 drout = 3.4946
+ pscbe1 = 4.5E8 pscbe2 = 1E-8 pvag = 0
+ delta = 0.01 fprout = 0 pdits = 1.4427E-15
+ pditsl = 0 pditsd = 0 lambda = 0
+ vtl = 0 lc = 0 xn = 0
+ alpha0 = 3.001670638882231E-4 lalpha0 = -3.608038759720174E-10 walpha0 = -1.783948583449416E-9
+ palpha0 = 3.637710787979964E-15 alpha1 = 0 beta0 = 15.827076836438899
+ lbeta0 = 1.070583336854855E-5 wbeta0 = -9.97696336801438E-6 pbeta0 = 2.042045900878358E-11
+ aigbacc = 1 bigbacc = 0 cigbacc = 0
+ nigbacc = 1 aigbinv = 0.35 bigbinv = 0.03
+ cigbinv = 6E-3 eigbinv = 1.1 nigbinv = 3
+ aigc = 0.43 bigc = 0.054 cigc = 0.075
+ aigsd = 0.43 bigsd = 0.054 cigsd = 0.075
+ dlcig = 0 nigc = 1 poxedge = 1
+ pigcd = 1 ntox = 1 toxref = 4.148E-9
+ agidl = 0 bgidl = 2.3E9 cgidl = 0.5
+ egidl = 0.8 noia = 9E41 noib = 1E27
+ noic = 8E11 em = 4.1E7 af = 1
+ ef = 1.2 kf = 0 lintnoi = -3E-7
+ tnoia = 2.5E7 tnoib = 9.9E6 ntnoi = 1
+ rnoia = 0.912 rnoib = 0.26 xpart = 0
+ cgso = {2.392894381E-10/sw_func_tox_lv_ratio} cgdo = {2.392894381E-10/sw_func_tox_lv_ratio} cgbo = {1E-14/sw_func_tox_lv_ratio}
+ ckappas = 0.6 cf = 1E-14 clc = 1E-7
+ cle = 0.6 dlc = 1.21071E-8 dwc = 2.6E-8
+ vfbcv = -1 noff = 3.8661 voffcv = -0.16994
+ acde = 0.38008 moin = 23.81 cgsl = {2.310725E-11/sw_func_tox_lv_ratio}
+ cgdl = {2.310725E-11/sw_func_tox_lv_ratio} ijthsrev = 0.1 ijthsfwd = 0.1
+ xjbvs = 1 bvs = 11.9 jss = 2.75E-3
+ jsws = 6E-10 cjs = {1.210E-03*sw_func_nsd_pw_cj} mjs = 0.42197
+ mjsws = 1E-3 cjsws = {3.230311424E-11*sw_func_nsd_pw_cj} cjswgs = {1.795291232E-10*sw_func_nsd_pw_cj}
+ mjswgs = 0.8 pbs = 0.7477 pbsws = 0.1
+ pbswgs = 0.79644 xrcrg1 = 12 xrcrg2 = 1
+ rbpb = 50 rbpd = 50 rbps = 50
+ rbdb = 50 rbsb = 50 gbmin = 1E-12
+ tnom = 30 ute = -0.55796572925 lute = -8.939266380284621E-7
+ wute = -2.983016510721E-6 pute = 3.713719208940679E-12 kt1 = -0.278545186337
+ lkt1 = 1.028580107335948E-7 wkt1 = 1.729725901664758E-7 pkt1 = -7.143845314653153E-13
+ kt1l = 0 kt2 = -0.0187382310889 lkt2 = -5.973551137198806E-8
+ wkt2 = -1.417074734247228E-7 pkt2 = 5.45173979872492E-13 ua1 = -5.973286598250007E-10
+ lua1 = 1.064936999713121E-14 wua1 = 1.88754961475241E-14 pua1 = -5.844043591523925E-20
+ ub1 = 5.124009045665005E-18 lub1 = -2.192491445117177E-23 wub1 = -4.349256327723045E-23
+ pub1 = 1.162124023728692E-28 uc1 = 2.264370932560003E-11 luc1 = -9.017788311661937E-17
+ wuc1 = -1.843193054867689E-16 puc1 = 2.028365909755966E-22 at = 1.931405051475551E6
+ lat = -3.748335456418715 wat = -9.171433079241528 pat = 1.835502342910561E-5
+ prt = 0 njs = 1.2928 xtis = 2
+ tpb = 1.2287E-3 tpbsw = 0 tpbswg = 0
+ tcj = 7.92E-4 tcjsw = 1E-5 tcjswg = 0
+ tvoff = 0 tvfbsdoff = 0 saref = 3E-6
+ sbref = 3E-6 wlod = 0 ku0 = -2.7E-8
+ kvsat = 0.2 kvth0 = 7.9E-9 tku0 = 0
+ llodku0 = 0 wlodku0 = 1 llodvth = 0
+ wlodvth = 1 lku0 = 0 wku0 = 0
+ pku0 = 0 lkvth0 = 0 wkvth0 = 3E-7
+ pkvth0 = 0 stk2 = 0 lodk2 = 1
+ steta0 = 0 lodeta0 = 1

.model nlowvt_model.12 nmos
+ level = 54 lmin = 1E-6 lmax = 2E-6 wmin = 5E-6
+ wmax = 7E-6 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 4.148E-9
+ toxm = 4.148E-9 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 9.999999999999999E22 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {2.6E-8+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {1.2025E-8-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = -1.33E-8 dwb = -1.08E-8 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = 0.449360133742969 lvth0 = -1.278750712539483E-8
+ wvth0 = -1.47368119017602E-7 pvth0 = 1.333637766056437E-13 vfb = 0
+ k1 = 0.120901197167 lk1 = 2.942707304878668E-7 wk1 = 2.140767132237686E-6
+ pk1 = -2.025700839467494E-12 k2 = 0.09714894945084 lk2 = -1.112971764322973E-7
+ wk2 = -7.740769182874964E-7 pk2 = 7.177564250829931E-13 k3 = 1.65
+ k3b = 1.6 w0 = 1E-7 lpe0 = 2.3802E-7
+ lpeb = -4.9152E-8 vbm = -3 dvtp0 = 0
+ dvtp1 = 0 dvt0 = 0.07665 dvt1 = 0.1252
+ dvt2 = -0.05637 dvt0w = 0 dvt1w = 5.3E6
+ dvt2w = -0.032 vfbsdoff = 0 u0 = 0.043068955775407
+ lu0 = -1.140052749945847E-8 wu0 = -3.354352848678794E-8 pu0 = 2.269640169816725E-14
+ ua = -8.808287691490269E-10 lua = -5.481909813836353E-16 wua = -4.815343405161107E-16
+ pua = 3.795197427777371E-23 ub = 2.774835794838001E-18 lub = 8.067765350985351E-26
+ wub = -1.091734198100431E-24 pub = 4.793263645671754E-31 uc = -7.966107077620006E-11
+ luc = 1.872781595380325E-16 wuc = 9.68039265288838E-16 puc = -1.118892262074714E-21
+ ud = 0 up = 0 lp = 1
+ eu = 1.67 vsat = 7.6405217763E3 lvsat = 0.05951408900862
+ wvsat = 0.080205947025268 pvsat = -5.234137826082753E-8 a0 = 2.49240933190194
+ la0 = -7.814814654764775E-7 wa0 = -2.097149036540918E-6 pa0 = 2.417840191304054E-12
+ ags = 0.872444940898898 lags = 1.563769800052621E-6 wags = -3.848322878077464E-7
+ pags = -1.817760709112745E-12 b0 = 0 b1 = 0
+ keta = 0.144161076744 lketa = -4.956360286513068E-7 wketa = -2.008508845863312E-6
+ pketa = 2.899825060327543E-12 a1 = 0 a2 = 0.38689047
+ rdsw = 103.65 rdswmin = 0 rdw = 0
+ rdwmin = 0 rsw = 0 rswmin = 0
+ prwb = 0 prwg = 0 wr = 1
+ voff = -0.141359674660307 lvoff = 2.809096347424863E-8 wvoff = 1.68777181680507E-7
+ pvoff = -1.790907162229198E-13 voffl = 0 minv = 0
+ nfactor = -0.173582824722337 lnfactor = 2.048641176403405E-6 wnfactor = 7.68951381924526E-6
+ pnfactor = -8.552554357587177E-12 eta0 = 7.506900318150001E-4 leta0 = -4.953509683648494E-10
+ weta0 = -1.10805137097462E-9 peta0 = 2.189454106477301E-15 etab = -5.873256246820002E-4
+ letab = 1.725510680903983E-10 wetab = 3.177364567185371E-10 petab = -6.278313516529934E-16
+ dsub = 0.175683046596022 ldsub = -4.6448472609231E-7 wdsub = -1.578677365703204E-6
+ pdsub = 7.819607662340774E-12 cit = 3.932225150000001E-5 lcit = -3.349680135142501E-11
+ wcit = -1.698265004220001E-10 pcit = 1.65742173086851E-16 cdsc = 3.8556E-37
+ cdscb = -1.1484E-4 cdscd = 4.7984E-6 pclm = 1.2154177404582
+ lpclm = -1.063127066020181E-6 wpclm = -6.852022662237577E-6 ppclm = 7.398531715989323E-12
+ pdiblc1 = 0.39 pdiblc2 = 0.01047271418283 lpdiblc2 = -3.968843342132936E-9
+ wpdiblc2 = -2.402207292280282E-8 ppdiblc2 = 5.058782606956861E-14 pdiblcb = 0
+ drout = 3.4946 pscbe1 = 4.5E8 pscbe2 = 1E-8
+ pvag = 0 delta = 0.01 fprout = 0
+ pdits = 1.4427E-15 pditsl = 0 pditsd = 0
+ lambda = 0 vtl = 0 lc = 0
+ xn = 0 alpha0 = 1.615313884173847E-4 lalpha0 = -8.686671302541434E-11
+ walpha0 = 1.741389270598548E-10 palpha0 = -2.31372228410829E-16 alpha1 = 0
+ beta0 = 20.70076232074269 lbeta0 = 1.075674535838471E-6 wbeta0 = 3.447517175213776E-6
+ pbeta0 = -6.105643320608098E-12 aigbacc = 1 bigbacc = 0
+ cigbacc = 0 nigbacc = 1 aigbinv = 0.35
+ bigbinv = 0.03 cigbinv = 6E-3 eigbinv = 1.1
+ nigbinv = 3 aigc = 0.43 bigc = 0.054
+ cigc = 0.075 aigsd = 0.43 bigsd = 0.054
+ cigsd = 0.075 dlcig = 0 nigc = 1
+ poxedge = 1 pigcd = 1 ntox = 1
+ toxref = 4.148E-9 agidl = 0 bgidl = 2.3E9
+ cgidl = 0.5 egidl = 0.8 noia = 9E41
+ noib = 1E27 noic = 8E11 em = 4.1E7
+ af = 1 ef = 1.2 kf = 0
+ lintnoi = -3E-7 tnoia = 2.5E7 tnoib = 9.9E6
+ ntnoi = 1 rnoia = 0.912 rnoib = 0.26
+ xpart = 0 cgso = {2.392894381E-10/sw_func_tox_lv_ratio} cgdo = {2.392894381E-10/sw_func_tox_lv_ratio}
+ cgbo = {1E-14/sw_func_tox_lv_ratio} ckappas = 0.6 cf = 1E-14
+ clc = 1E-7 cle = 0.6 dlc = 1.21071E-8
+ dwc = 2.6E-8 vfbcv = -1 noff = 3.8661
+ voffcv = -0.16994 acde = 0.38008 moin = 23.81
+ cgsl = {2.310725E-11/sw_func_tox_lv_ratio} cgdl = {2.310725E-11/sw_func_tox_lv_ratio} ijthsrev = 0.1
+ ijthsfwd = 0.1 xjbvs = 1 bvs = 11.9
+ jss = 2.75E-3 jsws = 6E-10 cjs = {1.210E-03*sw_func_nsd_pw_cj}
+ mjs = 0.42197 mjsws = 1E-3 cjsws = {3.230311424E-11*sw_func_nsd_pw_cj}
+ cjswgs = {1.795291232E-10*sw_func_nsd_pw_cj} mjswgs = 0.8 pbs = 0.7477
+ pbsws = 0.1 pbswgs = 0.79644 xrcrg1 = 12
+ xrcrg2 = 1 rbpb = 50 rbpd = 50
+ rbps = 50 rbdb = 50 rbsb = 50
+ gbmin = 1E-12 tnom = 30 ute = -1.40313207952
+ lute = 7.760798117875443E-7 wute = 5.4719689310496E-7 pute = -3.261805966349228E-12
+ kt1 = -0.21581645004 lkt1 = -2.109083575246185E-8 wkt1 = -2.422502253100794E-7
+ pkt1 = 1.06074990775584E-13 kt1l = 0 kt2 = -0.1388565097937
+ lkt2 = 1.776122014347615E-7 wkt2 = 6.455113927284277E-7 pkt2 = -1.010331138702826E-12
+ ua1 = 3.773859550759999E-9 lua1 = 2.01212065242578E-15 wua1 = -3.473293185240476E-15
+ pua1 = -1.428034563316309E-20 ub1 = -4.734467828669999E-18 lub1 = -2.445057071329518E-24
+ wub1 = 5.740125486599158E-24 pub1 = 1.893107100998013E-29 uc1 = 1.644089372665001E-10
+ luc1 = -3.702988852664408E-16 wuc1 = -1.063982251434042E-15 puc1 = 1.941006589020112E-21
+ at = 1.105105092299986E3 lat = 0.06584072263727 wat = 0.2076837456883
+ pat = -1.776424611144868E-7 prt = 0 njs = 1.2928
+ xtis = 2 tpb = 1.2287E-3 tpbsw = 0
+ tpbswg = 0 tcj = 7.92E-4 tcjsw = 1E-5
+ tcjswg = 0 tvoff = 0 tvfbsdoff = 0
+ saref = 3E-6 sbref = 3E-6 wlod = 0
+ ku0 = -2.7E-8 kvsat = 0.2 kvth0 = 7.9E-9
+ tku0 = 0 llodku0 = 0 wlodku0 = 1
+ llodvth = 0 wlodvth = 1 lku0 = 0
+ wku0 = 0 pku0 = 0 lkvth0 = 0
+ wkvth0 = 3E-7 pkvth0 = 0 stk2 = 0
+ lodk2 = 1 steta0 = 0 lodeta0 = 1

.model nlowvt_model.13 nmos
+ level = 54 lmin = 5E-7 lmax = 1E-6 wmin = 5E-6
+ wmax = 7E-6 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 4.148E-9
+ toxm = 4.148E-9 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 9.999999999999999E22 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {2.6E-8+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {1.2025E-8-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = -1.33E-8 dwb = -1.08E-8 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = 0.442438900423672 lvth0 = -6.032729467426532E-9
+ wvth0 = -6.236531162087886E-9 pvth0 = -4.373596561945227E-15 vfb = 0
+ k1 = 0.4491500363 lk1 = -2.608372406398503E-8 wk1 = -1.066590696924009E-7
+ pk1 = 1.67674762306174E-13 k2 = -0.019031533224547 lk2 = 2.089165634746849E-9
+ wk2 = 1.280933034282039E-8 pk2 = -5.020520926776456E-14 k3 = 1.65
+ k3b = 1.6 w0 = 1E-7 lpe0 = 2.3802E-7
+ lpeb = -4.9152E-8 vbm = -3 dvtp0 = 0
+ dvtp1 = 0 dvt0 = 0.07665 dvt1 = 0.1252
+ dvt2 = -0.05637 dvt0w = 0 dvt1w = 5.3E6
+ dvt2w = -0.032 vfbsdoff = 0 u0 = 0.0396199942462
+ lu0 = -8.034513495028899E-9 wu0 = -3.854594095151769E-8 pu0 = 2.757850614312026E-14
+ ua = -6.587525350002164E-10 lua = -7.64926282101167E-16 wua = -3.910682474857739E-15
+ pua = 3.384629095988486E-21 ub = 2.427710961534001E-18 lub = 4.194541345728923E-25
+ wub = 2.248286606349762E-24 pub = -2.78036693953599E-30 uc = 1.368390001917248E-10
+ luc = -2.401508472311381E-17 wuc = -2.043798722209041E-16 puc = 2.533019517791917E-23
+ ud = 0 up = 0 lp = 1
+ eu = 1.67 vsat = 1.458536264878801E5 lvsat = -0.075374990534647
+ wvsat = -0.891033466285471 pvsat = 8.955397271597876E-7 a0 = 2.165329138066441
+ la0 = -4.622675503027226E-7 wa0 = -1.005264539043949E-6 pa0 = 1.352215515971888E-12
+ ags = 0.556402918746401 lags = 1.872211011572352E-6 wags = 1.651645825230041E-5
+ pags = -1.83125752117313E-11 b0 = 0 b1 = 0
+ keta = -0.678927652109819 lketa = 3.076574162735776E-7 wketa = 1.726069439707383E-6
+ pketa = -7.449366174751766E-13 a1 = 0 a2 = 0.38689047
+ rdsw = 103.65 rdswmin = 0 rdw = 0
+ rdwmin = 0 rsw = 0 rswmin = 0
+ prwb = 0 prwg = 0 wr = 1
+ voff = -0.111021430915112 lvoff = -1.517645508874468E-9 wvoff = -2.743199372867014E-8
+ pvoff = 1.239962851766662E-14 voffl = 0 minv = 0
+ nfactor = 1.75811641390226 lnfactor = 1.633993044677296E-7 wnfactor = -2.85710442979702E-6
+ pnfactor = 1.740417722565634E-12 eta0 = 4.415009303699996E-4 leta0 = -1.935978648096013E-10
+ weta0 = 2.379728183637242E-9 peta0 = -1.214444349846145E-15 etab = -7.433104091044222E-4
+ letab = 3.247844184474608E-10 wetab = -6.252375366453537E-10 petab = 2.924641171704968E-16
+ dsub = -1.537953713533845 ldsub = 1.207939069956433E-6 wdsub = 1.255779497456547E-5
+ pdsub = -5.976882518144432E-12 cit = 5E-6 cdsc = 3.8556E-37
+ cdscb = -1.1484E-4 cdscd = 4.7984E-6 pclm = -0.557682842844
+ lpclm = 6.673304482536019E-7 wpclm = 3.588019492856114E-6 ppclm = -2.790427425274363E-12
+ pdiblc1 = 0.39 pdiblc2 = 1.003068750360001E-3 lpdiblc2 = 5.273057117686156E-9
+ wpdiblc2 = 6.461827838929872E-8 ppdiblc2 = -3.592072479347687E-14 pdiblcb = 0
+ drout = 3.4946 pscbe1 = 4.5E8 pscbe2 = 1E-8
+ pvag = 0 delta = 0.01 fprout = 0
+ pdits = 1.4427E-15 pditsl = 0 pditsd = 0
+ lambda = 0 vtl = 0 lc = 0
+ xn = 0 alpha0 = -1.048729175200697E-4 lalpha0 = 1.731305693542442E-10
+ walpha0 = 5.329990104004564E-10 palpha0 = -5.816017267470889E-16 alpha1 = 0
+ beta0 = 18.313320589144002 lbeta0 = 3.405698293792213E-6 wbeta0 = 1.719912311525066E-6
+ pbeta0 = -4.419587353891102E-12 aigbacc = 1 bigbacc = 0
+ cigbacc = 0 nigbacc = 1 aigbinv = 0.35
+ bigbinv = 0.03 cigbinv = 6E-3 eigbinv = 1.1
+ nigbinv = 3 aigc = 0.43 bigc = 0.054
+ cigc = 0.075 aigsd = 0.43 bigsd = 0.054
+ cigsd = 0.075 dlcig = 0 nigc = 1
+ poxedge = 1 pigcd = 1 ntox = 1
+ toxref = 4.148E-9 agidl = 0 bgidl = 2.3E9
+ cgidl = 0.5 egidl = 0.8 noia = 9E41
+ noib = 1E27 noic = 8E11 em = 4.1E7
+ af = 1 ef = 1.2 kf = 0
+ lintnoi = -3E-7 tnoia = 2.5E7 tnoib = 9.9E6
+ ntnoi = 1 rnoia = 0.912 rnoib = 0.26
+ xpart = 0 cgso = {2.392894381E-10/sw_func_tox_lv_ratio} cgdo = {2.392894381E-10/sw_func_tox_lv_ratio}
+ cgbo = {1E-14/sw_func_tox_lv_ratio} ckappas = 0.6 cf = 1E-14
+ clc = 1E-7 cle = 0.6 dlc = 1.21071E-8
+ dwc = 2.6E-8 vfbcv = -1 noff = 3.8661
+ voffcv = -0.16994 acde = 0.38008 moin = 23.81
+ cgsl = {2.310725E-11/sw_func_tox_lv_ratio} cgdl = {2.310725E-11/sw_func_tox_lv_ratio} ijthsrev = 0.1
+ ijthsfwd = 0.1 xjbvs = 1 bvs = 11.9
+ jss = 2.75E-3 jsws = 6E-10 cjs = {1.210E-03*sw_func_nsd_pw_cj}
+ mjs = 0.42197 mjsws = 1E-3 cjsws = {3.230311424E-11*sw_func_nsd_pw_cj}
+ cjswgs = {1.795291232E-10*sw_func_nsd_pw_cj} mjswgs = 0.8 pbs = 0.7477
+ pbsws = 0.1 pbswgs = 0.79644 xrcrg1 = 12
+ xrcrg2 = 1 rbpb = 50 rbpd = 50
+ rbps = 50 rbdb = 50 rbsb = 50
+ gbmin = 1E-12 tnom = 30 ute = -0.288159259839999
+ lute = -3.120779115791525E-7 wute = -4.981024536151685E-6 pute = 2.133461737533795E-12
+ kt1 = -0.219377453922 lkt1 = -1.761547401382403E-8 wkt1 = -2.175011166259435E-7
+ pkt1 = 8.192109815530155E-14 kt1l = 0 kt2 = 0.0863442531484
+ lkt2 = -4.217248315858099E-8 wkt2 = -6.092041560242836E-7 pkt2 = 2.142085011023825E-13
+ ua1 = 9.152284981160002E-9 lua1 = -3.236953646373103E-15 wua1 = -3.55905591603797E-14
+ pua1 = 1.706450009527404E-20 ub1 = -1.18674032778E-17 lub1 = 4.516331280248913E-24
+ wub1 = 4.989423769219443E-23 pub1 = -2.416113479707058E-29 uc1 = -5.094243914242403E-10
+ luc1 = 2.873287518692872E-16 wuc1 = 2.371965846314341E-15 puc1 = -1.412306956977423E-21
+ at = 1.360319227019999E4 lat = 0.053643214455998 wat = 0.40826907283505
+ pat = -3.734037111433583E-7 prt = 0 njs = 1.2928
+ xtis = 2 tpb = 1.2287E-3 tpbsw = 0
+ tpbswg = 0 tcj = 7.92E-4 tcjsw = 1E-5
+ tcjswg = 0 tvoff = 0 tvfbsdoff = 0
+ saref = 2.74E-6 sbref = 2.74E-6 wlod = 0
+ ku0 = -2.7E-8 kvsat = 0.2 kvth0 = 7.9E-9
+ tku0 = 0 llodku0 = 0 wlodku0 = 1
+ llodvth = 0 wlodvth = 1 lku0 = 0
+ wku0 = 0 pku0 = 0 lkvth0 = 0
+ wkvth0 = 3E-7 pkvth0 = 0 stk2 = 0
+ lodk2 = 1 steta0 = 0 lodeta0 = 1

.model nlowvt_model.14 nmos
+ level = 54 lmin = 2.5E-7 lmax = 5E-7 wmin = 5E-6
+ wmax = 7E-6 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 4.148E-9
+ toxm = 4.148E-9 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 9.999999999999999E22 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {2.6E-8+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {1.2025E-8-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = -1.33E-8 dwb = -1.08E-8 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = 0.49409312589808 lvth0 = -3.06175580819712E-8
+ wvth0 = 1.023309765037895E-8 pvth0 = -1.221231639523882E-14 vfb = 0
+ k1 = 0.274337228448 lk1 = 5.711843183317426E-8 wk1 = 1.362642562632939E-7
+ pk1 = 5.205540531756104E-14 k2 = 0.025328257138548 lk2 = -1.90238765885683E-8
+ wk2 = -7.788159514699783E-8 pk2 = -7.040863280885588E-15 k3 = 1.65
+ k3b = 1.6 w0 = 1E-7 lpe0 = 2.3802E-7
+ lpeb = -4.9152E-8 vbm = -3 dvtp0 = 0
+ dvtp1 = 0 dvt0 = 0.07665 dvt1 = 0.1252
+ dvt2 = -0.05637 dvt0w = 0 dvt1w = 5.3E6
+ dvt2w = -0.032 vfbsdoff = 0 u0 = 0.026667460588592
+ lu0 = -1.86975510069036E-9 wu0 = 8.256575060126837E-9 pu0 = 5.302848647378043E-15
+ ua = -2.009938431041719E-9 lua = -1.218293548802136E-16 wua = 2.253231119670908E-15
+ pua = 4.509144206725761E-22 ub = 3.202014313104001E-18 lub = 5.092445439315084E-26
+ wub = -2.675582732774599E-24 pub = -4.368513275797508E-31 uc = 1.326514729124885E-10
+ luc = -2.202203111456128E-17 wuc = -4.078240413127947E-16 puc = 1.221594474572045E-22
+ ud = 0 up = 0 lp = 1
+ eu = 1.67 vsat = -1.883775500551482E5 lvsat = 0.083702337941008
+ wvsat = 1.994070018836074 pvsat = -4.776252765838113E-7 a0 = 0.442084651559999
+ la0 = 3.579106630500181E-7 wa0 = 6.087953829201124E-6 pa0 = -2.023801766394354E-12
+ ags = 8.548123922998805 lags = -1.931448600401579E-6 wags = -4.180626762619568E-5
+ pags = 9.446126170138912E-12 b0 = 0 b1 = 0
+ keta = -0.126459204411073 lketa = 4.471005859135964E-8 wketa = 7.839564433150359E-7
+ pketa = -2.965379368422388E-13 a1 = 0 a2 = 0.38689047
+ rdsw = 103.65 rdswmin = 0 rdw = 0
+ rdwmin = 0 rsw = 0 rswmin = 0
+ prwb = 0 prwg = 0 wr = 1
+ voff = -0.123016791094264 lvoff = 4.191546168392951E-9 wvoff = 3.039438128086632E-8
+ pvoff = -1.512283466812225E-14 voffl = 0 minv = 0
+ nfactor = 1.8237772575086 lnfactor = 1.321480259532918E-7 wnfactor = 1.116696043923844E-6
+ pnfactor = -1.509126129018104E-13 eta0 = -0.010040261618129 leta0 = 4.795197020148708E-9
+ weta0 = 3.364616062520793E-8 peta0 = -1.609570287041171E-14 etab = -0.040163080603906
+ letab = 1.908662404266306E-8 wetab = 4.496645557569889E-7 petab = -2.140229630009347E-13
+ dsub = 1.814680033366508 ldsub = -3.877469618807893E-7 wdsub = -1.077280427338129E-6
+ pdsub = 5.127316193915823E-13 cit = 5E-6 cdsc = 3.8556E-37
+ cdscb = -1.1484E-4 cdscd = 4.7984E-6 pclm = 1.291626919616
+ lpclm = -2.128485331892352E-7 wpclm = -4.522549177003969E-6 ppclm = 1.069797733145543E-12
+ pdiblc1 = 0.39 pdiblc2 = 0.01258209612768 lpdiblc2 = -2.379809625492954E-10
+ wpdiblc2 = -3.580996370552063E-8 ppdiblc2 = 1.187809703155239E-14 pdiblcb = 0
+ drout = 3.4946 pscbe1 = 4.5E8 pscbe2 = 1E-8
+ pvag = 0 delta = 0.01 fprout = 0
+ pdits = 1.4427E-15 pditsl = 0 pditsd = 0
+ lambda = 0 vtl = 0 lc = 0
+ xn = 0 alpha0 = -4.373541746579454E-3 lalpha0 = 2.204803498545058E-9
+ walpha0 = 1.452184349430479E-8 palpha0 = -7.239592258861357E-15 alpha1 = 0
+ beta0 = 18.502665043792398 lbeta0 = 3.315579800602307E-6 wbeta0 = -2.420894062020003E-6
+ pbeta0 = -2.448770560402326E-12 aigbacc = 1 bigbacc = 0
+ cigbacc = 0 nigbacc = 1 aigbinv = 0.35
+ bigbinv = 0.03 cigbinv = 6E-3 eigbinv = 1.1
+ nigbinv = 3 aigc = 0.43 bigc = 0.054
+ cigc = 0.075 aigsd = 0.43 bigsd = 0.054
+ cigsd = 0.075 dlcig = 0 nigc = 1
+ poxedge = 1 pigcd = 1 ntox = 1
+ toxref = 4.148E-9 agidl = 0 bgidl = 2.3E9
+ cgidl = 0.5 egidl = 0.8 noia = 9E41
+ noib = 1E27 noic = 8E11 em = 4.1E7
+ af = 1 ef = 1.2 kf = 0
+ lintnoi = -3E-7 tnoia = 2.5E7 tnoib = 9.9E6
+ ntnoi = 1 rnoia = 0.912 rnoib = 0.26
+ xpart = 0 cgso = {2.392894381E-10/sw_func_tox_lv_ratio} cgdo = {2.392894381E-10/sw_func_tox_lv_ratio}
+ cgbo = {1E-14/sw_func_tox_lv_ratio} ckappas = 0.6 cf = 1E-14
+ clc = 1E-7 cle = 0.6 dlc = 1.21071E-8
+ dwc = 2.6E-8 vfbcv = -1 noff = 3.8661
+ voffcv = -0.16994 acde = 0.38008 moin = 23.81
+ cgsl = {2.310725E-11/sw_func_tox_lv_ratio} cgdl = {2.310725E-11/sw_func_tox_lv_ratio} ijthsrev = 0.1
+ ijthsfwd = 0.1 xjbvs = 1 bvs = 11.9
+ jss = 2.75E-3 jsws = 6E-10 cjs = {1.210E-03*sw_func_nsd_pw_cj}
+ mjs = 0.42197 mjsws = 1E-3 cjsws = {3.230311424E-11*sw_func_nsd_pw_cj}
+ cjswgs = {1.795291232E-10*sw_func_nsd_pw_cj} mjswgs = 0.8 pbs = 0.7477
+ pbsws = 0.1 pbswgs = 0.79644 xrcrg1 = 12
+ xrcrg2 = 1 rbpb = 50 rbpd = 50
+ rbps = 50 rbdb = 50 rbsb = 50
+ gbmin = 1E-12 tnom = 30 ute = 1.560464487992001
+ lute = -1.191930384359793E-6 wute = -1.380733509896842E-5 pute = 6.334344249906419E-12
+ kt1 = -0.180713990204 lkt1 = -3.601734957040623E-8 wkt1 = -5.088109042306091E-7
+ pkt1 = 2.205699915657421E-13 kt1l = 0 kt2 = 5.646006553200024E-3
+ lkt2 = -3.764152691595543E-9 wkt2 = -2.362118087868337E-7 pkt2 = 3.668279343471826E-14
+ ua1 = 8.609815863764002E-9 lua1 = -2.978765469948476E-15 wua1 = -3.129738521214428E-14
+ pua1 = 1.502116395461139E-20 ub1 = -7.617292603724E-18 lub1 = 2.493491104922438E-24
+ wub1 = 2.421685975466636E-23 pub1 = -1.193998676770409E-29 uc1 = 2.941949073292801E-10
+ luc1 = -9.515385337245082E-17 wuc1 = -1.701123983999678E-15 puc1 = 5.262801477605345E-22
+ at = 1.759026985984E5 lat = -0.023603235580908 wat = -0.614468824808084
+ pat = 1.133683912398912E-7 prt = 0 njs = 1.2928
+ xtis = 2 tpb = 1.2287E-3 tpbsw = 0
+ tpbswg = 0 tcj = 7.92E-4 tcjsw = 1E-5
+ tcjswg = 0 tvoff = 0 tvfbsdoff = 0
+ saref = 1.74E-6 sbref = 1.74E-6 wlod = 0
+ ku0 = -2.7E-8 kvsat = 0.2 kvth0 = 7.9E-9
+ tku0 = 0 llodku0 = 0 wlodku0 = 1
+ llodvth = 0 wlodvth = 1 lku0 = 0
+ wku0 = 0 pku0 = 0 lkvth0 = 0
+ wkvth0 = 3E-7 pkvth0 = 0 stk2 = 0
+ lodk2 = 1 steta0 = 0 lodeta0 = 1

.model nlowvt_model.15 nmos
+ level = 54 lmin = 1.8E-7 lmax = 2.5E-7 wmin = 5E-6
+ wmax = 7E-6 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 4.148E-9
+ toxm = 4.148E-9 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 9.999999999999999E22 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {2.6E-8+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {1.2025E-8-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = -1.33E-8 dwb = -1.08E-8 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = 0.648283385811429 lvth0 = -6.545684730939229E-8
+ wvth0 = -2.75732725609235E-7 pvth0 = 5.240166137027096E-14 vfb = 0
+ k1 = 0.173405973299999 lk1 = 7.992384893386513E-8 wk1 = 9.881835550544618E-7
+ pk1 = -1.404357602443033E-13 k2 = 0.035285514399037 lk2 = -2.127371886657584E-8
+ wk2 = -2.751469173797617E-7 pk2 = 3.75312362776074E-14 k3 = 1.65
+ k3b = 1.6 w0 = 1E-7 lpe0 = 2.3802E-7
+ lpeb = -4.9152E-8 vbm = -3 dvtp0 = 0
+ dvtp1 = 0 dvt0 = 0.07665 dvt1 = 0.1252
+ dvt2 = -0.05637 dvt0w = 0 dvt1w = 5.3E6
+ dvt2w = -0.032 vfbsdoff = 0 u0 = 0.021625997380114
+ lu0 = -7.306364887348211E-10 wu0 = 1.23161377535566E-7 pu0 = -2.065989147194743E-14
+ ua = -3.118749799151573E-9 lua = 1.28706573744208E-16 wua = 1.517871540335028E-14
+ pua = -2.469598753224776E-21 ub = 4.650873680085714E-18 lub = -2.764453195763671E-25
+ wub = -1.42218974393784E-23 pub = 2.172038480377378E-30 uc = -9.41980474406435E-12
+ luc = 1.007897407193683E-17 wuc = 6.434596423904192E-16 puc = -1.153781008755367E-22
+ ud = 0 up = 0 lp = 1
+ eu = 1.67 vsat = 2.005434251085285E5 lvsat = -4.174356397225023E-3
+ wvsat = -0.336420639092428 pvsat = 4.894908757513347E-8 a0 = 6.539995572428571
+ la0 = -1.019912309520236E-6 wa0 = -9.260408552662292E-6 pa0 = 1.444160713787684E-12
+ ags = -2.747483879571429 lags = 6.207939825891643E-7 wags = 4.55715505548001E-7
+ pags = -1.029689184785708E-13 b0 = 0 b1 = 0
+ keta = 0.67324190717929 lketa = -1.359824075724828E-7 wketa = -2.965922873327819E-6
+ pketa = 5.507472947532142E-13 a1 = 0 a2 = 0.38689047
+ rdsw = 103.65 rdswmin = 0 rdw = 0
+ rdwmin = 0 rsw = 0 rswmin = 0
+ prwb = 0 prwg = 0 wr = 1
+ voff = -0.174140511097401 lvoff = 1.574295070310184E-8 wvoff = 7.086108771418797E-8
+ pvoff = -2.426628698673128E-14 voffl = 0 minv = 0
+ nfactor = 1.258837744743143 lnfactor = 2.597961088626469E-7 wnfactor = -5.070913600364264E-8
+ pnfactor = 1.128625875028051E-13 eta0 = -0.061889163338682 leta0 = 1.651045636390755E-8
+ weta0 = -6.392919289844428E-7 peta0 = 1.359546584768888E-13 etab = 0.164131862569436
+ letab = -2.70738183673534E-8 wetab = -1.523151754861823E-6 petab = 2.317348823833857E-13
+ dsub = -0.420490721224671 ldsub = 1.172898701190875E-7 wdsub = 3.997624737363845E-6
+ pdsub = -6.339432025728283E-13 cit = -4.254565381657653E-8 lcit = 1.139363190479856E-12
+ wcit = 3.503560720271758E-11 pcit = -7.916295447454037E-18 cdsc = 3.8556E-37
+ cdscb = -1.1484E-4 cdscd = 4.7984E-6 pclm = 0.736800603785714
+ lpclm = -8.748552712738207E-8 wpclm = 1.110144217554002E-6 ppclm = -2.029093393548306E-13
+ pdiblc1 = -0.969000904251971 lpdiblc1 = 3.070662543157329E-7 wpdiblc1 = 5.591131412638944E-11
+ ppdiblc1 = -1.263316142685769E-17 pdiblc2 = -0.013008331911429 lpdiblc2 = 5.544176252887287E-9
+ wpdiblc2 = 1.908506004034629E-7 ppdiblc2 = -3.933585742887244E-14 pdiblcb = 0
+ drout = 3.4946 pscbe1 = 4.5E8 pscbe2 = 1E-8
+ pvag = 0 delta = 0.01 fprout = 0
+ pdits = 1.4427E-15 pditsl = 0 pditsd = 0
+ lambda = 0 vtl = 0 lc = 0
+ xn = 0 alpha0 = 0.020529807773742 lalpha0 = -3.422108325571543E-9
+ walpha0 = -8.839497358119219E-8 palpha0 = 1.601446255934718E-14 alpha1 = 0
+ beta0 = 50.14962747264711 lbeta0 = -3.835051360197413E-6 wbeta0 = -9.605904176188931E-5
+ pbeta0 = 1.870876891238314E-11 aigbacc = 1 bigbacc = 0
+ cigbacc = 0 nigbacc = 1 aigbinv = 0.35
+ bigbinv = 0.03 cigbinv = 6E-3 eigbinv = 1.1
+ nigbinv = 3 aigc = 0.43 bigc = 0.054
+ cigc = 0.075 aigsd = 0.43 bigsd = 0.054
+ cigsd = 0.075 dlcig = 0 nigc = 1
+ poxedge = 1 pigcd = 1 ntox = 1
+ toxref = 4.148E-9 agidl = 0 bgidl = 2.3E9
+ cgidl = 0.5 egidl = 0.8 noia = 9E41
+ noib = 1E27 noic = 8E11 em = 4.1E7
+ af = 1 ef = 1.2 kf = 0
+ lintnoi = -3E-7 tnoia = 2.5E7 tnoib = 9.9E6
+ ntnoi = 1 rnoia = 0.912 rnoib = 0.26
+ xpart = 0 cgso = {2.392894381E-10/sw_func_tox_lv_ratio} cgdo = {2.392894381E-10/sw_func_tox_lv_ratio}
+ cgbo = {1E-14/sw_func_tox_lv_ratio} ckappas = 0.6 cf = 1E-14
+ clc = 1E-7 cle = 0.6 dlc = 1.21071E-8
+ dwc = 2.6E-8 vfbcv = -1 noff = 3.8661
+ voffcv = -0.16994 acde = 0.38008 moin = 23.81
+ cgsl = {2.310725E-11/sw_func_tox_lv_ratio} cgdl = {2.310725E-11/sw_func_tox_lv_ratio} ijthsrev = 0.1
+ ijthsfwd = 0.1 xjbvs = 1 bvs = 11.9
+ jss = 2.75E-3 jsws = 6E-10 cjs = {1.210E-03*sw_func_nsd_pw_cj}
+ mjs = 0.42197 mjsws = 1E-3 cjsws = {3.230311424E-11*sw_func_nsd_pw_cj}
+ cjswgs = {1.795291232E-10*sw_func_nsd_pw_cj} mjswgs = 0.8 pbs = 0.7477
+ pbsws = 0.1 pbswgs = 0.79644 xrcrg1 = 12
+ xrcrg2 = 1 rbpb = 50 rbpd = 50
+ rbps = 50 rbdb = 50 rbsb = 50
+ gbmin = 1E-12 tnom = 30 ute = -6.012811911400004
+ lute = 5.192514180828304E-7 wute = 3.385946941869293E-5 pute = -4.435970230859162E-12
+ kt1 = -0.374009114 lkt1 = 7.657683651300014E-9 wkt1 = 1.332854987214858E-6
+ pkt1 = -1.955544166063611E-13 kt1l = 0 kt2 = -0.086782857302857
+ lkt2 = 1.712014909668058E-8 wkt2 = 3.59028789305966E-7 pkt2 = -9.78118197043498E-14
+ ua1 = -1.33158405701943E-8 lua1 = 1.9753366013044E-15 wua1 = 1.0323024246315E-13
+ pua1 = -1.537535351862134E-20 ub1 = 1.103545863191429E-17 lub1 = -1.721098036770034E-24
+ wub1 = -9.05419013133405E-23 pub1 = 1.398975529561205E-29 uc1 = -4.242991203064288E-10
+ luc1 = 6.718987217183756E-17 wuc1 = 2.09943204727621E-15 puc1 = -3.324554875062522E-22
+ at = 6.959335782E4 lat = 4.173599679709964E-4 wat = -0.482584942901932
+ pat = 8.356922812319624E-8 prt = 0 njs = 1.2928
+ xtis = 2 tpb = 1.2287E-3 tpbsw = 0
+ tpbswg = 0 tcj = 7.92E-4 tcjsw = 1E-5
+ tcjswg = 0 tvoff = 0 tvfbsdoff = 0
+ saref = 1.25E-6 sbref = 1.24E-6 wlod = 0
+ ku0 = -2.7E-8 kvsat = 0.2 kvth0 = 7.9E-9
+ tku0 = 0 llodku0 = 0 wlodku0 = 1
+ llodvth = 0 wlodvth = 1 lku0 = 0
+ wku0 = 0 pku0 = 0 lkvth0 = 0
+ wkvth0 = 3E-7 pkvth0 = 0 stk2 = 0
+ lodk2 = 1 steta0 = 0 lodeta0 = 1

.model nlowvt_model.16 nmos
+ level = 54 lmin = 1.5E-7 lmax = 1.8E-7 wmin = 5E-6
+ wmax = 7E-6 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 4.148E-9
+ toxm = 4.148E-9 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 9.999999999999999E22 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {2.6E-8+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {1.2025E-8-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = -1.33E-8 dwb = -1.08E-8 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = 0.239953534053333 lvth0 = -1.777806927717355E-9
+ wvth0 = 6.952038603743944E-8 pvth0 = -1.440561391027848E-15 vfb = 0
+ k1 = 1.569238482733334 lk1 = -1.377562309122634E-7 wk1 = -3.877168928431202E-6
+ pk1 = 6.183159595552858E-13 k2 = -0.383875840304047 lk2 = 4.40944943993701E-8
+ wk2 = 1.156822877603556E-6 pk2 = -1.85784453250041E-13 k3 = 1.65
+ k3b = 1.6 w0 = 1E-7 lpe0 = 2.3802E-7
+ lpeb = -4.9152E-8 vbm = -3 dvtp0 = 0
+ dvtp1 = 0 dvt0 = 0.07665 dvt1 = 0.1252
+ dvt2 = -0.05637 dvt0w = 0 dvt1w = 5.3E6
+ dvt2w = -0.032 vfbsdoff = 0 u0 = 0.0194266354008
+ lu0 = -3.876459880607626E-10 wu0 = -3.624021112335854E-8 pu0 = 4.198786279411848E-15
+ ua = -6.754774968259666E-9 lua = 6.95744698866615E-16 wua = 2.263605105662217E-14
+ pua = -3.632570248352528E-21 ub = 1.013281276256667E-17 lub = -1.131353719489272E-24
+ wub = -3.858500174851322E-23 pub = 5.971464597386952E-30 uc = 4.022738493443334E-10
+ luc = -5.412465128314879E-17 wuc = -1.500101023342429E-15 puc = 2.189101849455009E-22
+ ud = 0 up = 0 lp = 1
+ eu = 1.67 vsat = 1.519079454683002E5 lvsat = 3.410346652668585E-3
+ wvsat = 0.208978980550851 pvsat = -3.610598310823574E-8 a0 = 0
+ ags = 1.165531559333332 lags = 1.055922489196682E-8 wags = -1.113852820247997E-6
+ pags = 1.41805261929315E-13 b0 = 0 b1 = 0
+ keta = 0.580818027040581 lketa = -1.215689034648511E-7 wketa = -2.945183695305553E-6
+ pketa = 5.475130199406418E-13 a1 = 0 a2 = 0.38689047
+ rdsw = 103.65 rdswmin = 0 rdw = 0
+ rdwmin = 0 rsw = 0 rswmin = 0
+ prwb = 0 prwg = 0 wr = 1
+ voff = -0.40861810149534 lvoff = 5.23097309256604E-8 wvoff = 2.009846450931504E-6
+ pvoff = -3.266510543804716E-13 voffl = 0 minv = 0
+ nfactor = -3.821753976047002 lnfactor = 1.05211438771987E-6 wnfactor = 3.158014253793255E-5
+ pnfactor = -4.819968731047545E-12 eta0 = -0.298021796609047 leta0 = 5.333534052242097E-8
+ weta0 = 2.540599762844978E-6 peta0 = -3.599494508639093E-13 etab = -0.172255637842827
+ letab = 2.538581232193893E-8 wetab = 6.612992731958603E-7 petab = -1.089302554422099E-13
+ dsub = 0.632244738136666 ldsub = -4.688422476831312E-8 wdsub = -3.504541593645585E-7
+ pdsub = 4.413970137196614E-14 cit = 1.676593985890536E-5 lcit = -1.481920125229129E-12
+ wcit = -8.174975013967436E-11 pcit = 1.029638103009198E-17 cdsc = 3.8556E-37
+ cdscb = -1.1484E-4 cdscd = 4.7984E-6 pclm = 1.325293189233334
+ lpclm = -1.792609458279384E-7 wpclm = -8.604881031793201E-6 ppclm = 1.312148848280866E-12
+ pdiblc1 = 8.805549376714167 lpdiblc1 = -1.217274862000936E-6 wpdiblc1 = -3.628149135934864E-5
+ ppdiblc1 = 5.658094663698432E-12 pdiblc2 = 0.124956462306333 lpdiblc2 = -1.597143340537269E-8
+ wpdiblc2 = -4.184131420184043E-7 ppdiblc2 = 5.567882320181773E-14 pdiblcb = 0
+ drout = 3.4946 pscbe1 = 4.5E8 pscbe2 = 1E-8
+ pvag = 0 delta = 0.01 fprout = 0
+ pdits = 1.4427E-15 pditsl = 0 pditsd = 0
+ lambda = 0 vtl = 0 lc = 0
+ xn = 0 alpha0 = -6.393844807937837E-3 lalpha0 = 7.766352945414054E-10
+ walpha0 = 5.614854197816409E-8 palpha0 = -6.527098692134426E-15 alpha1 = 0
+ beta0 = 20.667706561966668 lbeta0 = 7.62654205823198E-7 wbeta0 = 7.346207433913558E-5
+ pbeta0 = -7.728049143571676E-12 aigbacc = 1 bigbacc = 0
+ cigbacc = 0 nigbacc = 1 aigbinv = 0.35
+ bigbinv = 0.03 cigbinv = 6E-3 eigbinv = 1.1
+ nigbinv = 3 aigc = 0.43 bigc = 0.054
+ cigc = 0.075 aigsd = 0.43 bigsd = 0.054
+ cigsd = 0.075 dlcig = 0 nigc = 1
+ poxedge = 1 pigcd = 1 ntox = 1
+ toxref = 4.148E-9 agidl = 0 bgidl = 2.3E9
+ cgidl = 0.5 egidl = 0.8 noia = 9E41
+ noib = 1E27 noic = 8E11 em = 4.1E7
+ af = 1 ef = 1.2 kf = 0
+ lintnoi = -3E-7 tnoia = 2.5E7 tnoib = 9.9E6
+ ntnoi = 1 rnoia = 0.912 rnoib = 0.26
+ xpart = 0 cgso = {2.392894381E-10/sw_func_tox_lv_ratio} cgdo = {2.392894381E-10/sw_func_tox_lv_ratio}
+ cgbo = {1E-14/sw_func_tox_lv_ratio} ckappas = 0.6 cf = 1E-14
+ clc = 1E-7 cle = 0.6 dlc = 1.21071E-8
+ dwc = 2.6E-8 vfbcv = -1 noff = 3.8661
+ voffcv = -0.16994 acde = 0.38008 moin = 23.81
+ cgsl = {2.310725E-11/sw_func_tox_lv_ratio} cgdl = {2.310725E-11/sw_func_tox_lv_ratio} ijthsrev = 0.1
+ ijthsfwd = 0.1 xjbvs = 1 bvs = 11.9
+ jss = 2.75E-3 jsws = 6E-10 cjs = {1.210E-03*sw_func_nsd_pw_cj}
+ mjs = 0.42197 mjsws = 1E-3 cjsws = {3.230311424E-11*sw_func_nsd_pw_cj}
+ cjswgs = {1.795291232E-10*sw_func_nsd_pw_cj} mjswgs = 0.8 pbs = 0.7477
+ pbsws = 0.1 pbswgs = 0.79644 xrcrg1 = 12
+ xrcrg2 = 1 rbpb = 50 rbpd = 50
+ rbps = 50 rbdb = 50 rbsb = 50
+ gbmin = 1E-12 tnom = 30 ute = -4.228318418333331
+ lute = 2.409596578390829E-7 wute = 9.636393704579987E-6 pute = -6.583815732432488E-13
+ kt1 = 0.078247527066667 lkt1 = -6.287173952304674E-8 wkt1 = -2.594152830259203E-6
+ pkt1 = 4.168624525287186E-13 kt1l = 0 kt2 = 0.350932040936667
+ lkt2 = -5.114148928377321E-8 wkt2 = -2.290785204987961E-6 pkt2 = 3.154266727057882E-13
+ ua1 = -6.71898347614667E-9 lua1 = 9.46556737487673E-16 wua1 = 2.980665184990706E-14
+ pua1 = -3.92494456248611E-21 ub1 = 5.84802748786667E-18 lub1 = -9.12118149855807E-25
+ wub1 = -2.364854552489761E-23 pub1 = 3.557736460404386E-30 uc1 = -2.500259603916669E-10
+ luc1 = 4.001197288313045E-17 wuc1 = 1.773413341671301E-15 puc1 = -2.816128703671668E-22
+ at = -7.223001372000013E4 lat = 0.022534714759634 wat = 0.946132531126561
+ pat = -1.392392619515471E-7 prt = 0 njs = 1.2928
+ xtis = 2 tpb = 1.2287E-3 tpbsw = 0
+ tpbswg = 0 tcj = 7.92E-4 tcjsw = 1E-5
+ tcjswg = 0 tvoff = 0 tvfbsdoff = 0
+ saref = 1.1E-6 sbref = 1.1E-6 wlod = 0
+ ku0 = -2.7E-8 kvsat = 0.2 kvth0 = 7.9E-9
+ tku0 = 0 llodku0 = 0 wlodku0 = 1
+ llodvth = 0 wlodvth = 1 lku0 = 0
+ wku0 = 0 pku0 = 0 lkvth0 = 0
+ wkvth0 = 3E-7 pkvth0 = 0 stk2 = 0
+ lodk2 = 1 steta0 = 0 lodeta0 = 1

.model nlowvt_model.17 nmos
+ level = 54 lmin = 8E-6 lmax = 2.02E-5 wmin = 3E-6
+ wmax = 5E-6 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 4.148E-9
+ toxm = 4.148E-9 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 9.999999999999999E22 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {2.6E-8+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {1.2025E-8-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = -1.33E-8 dwb = -1.08E-8 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = 0.428625 vfb = 0
+ k1 = 0.24736776 wk1 = 7.567582035200001E-7 k2 = 0.05125898698
+ wk2 = -2.958932598450399E-7 k3 = 1.65 k3b = 1.6
+ w0 = 1E-7 lpe0 = 2.3802E-7 lpeb = -4.9152E-8
+ vbm = -3 dvtp0 = 0 dvtp1 = 0
+ dvt0 = 0.07665 dvt1 = 0.1252 dvt2 = -0.05637
+ dvt0w = 0 dvt1w = 5.3E6 dvt2w = -0.032
+ vfbsdoff = 0 u0 = 0.0320233044 wu0 = 1.855428748799963E-9
+ ua = -1.508486209E-9 wua = 1.201240601131999E-15 ub = 2.94084734E-18
+ wub = -1.385080478320001E-24 uc = 7.254987096200001E-11 wuc = -1.043469351997604E-17
+ ud = 0 up = 0 lp = 1
+ eu = 1.67 vsat = 3.5078784E5 wvsat = -0.53358163232
+ a0 = 2.2794517696 wa0 = -1.754929275580798E-6 ags = 0.565636564
+ wags = -8.960612267200013E-8 b0 = 0 b1 = 0
+ keta = 0 a1 = 0 a2 = 0.38689047
+ rdsw = 103.65 rdswmin = 0 rdw = 0
+ rdwmin = 0 rsw = 0 rswmin = 0
+ prwb = 0 prwg = 0 wr = 1
+ voff = -0.1249454834 wvoff = 2.989617918319996E-8 voffl = 0
+ minv = 0 nfactor = 0.5601947258 wnfactor = 2.282660910261599E-6
+ eta0 = 0.08 etab = -0.07 dsub = 0.56
+ cit = 1.737E-5 wcit = -3.646676E-11 cdsc = 3.8556E-37
+ cdscb = -1.1484E-4 cdscd = 4.7984E-6 pclm = -0.125464596
+ wpclm = 9.59469629008E-7 pdiblc1 = 0.39 pdiblc2 = 6.403487E-3
+ wpdiblc2 = 9.08022323999997E-10 pdiblcb = 0 drout = 3.4946
+ pscbe1 = 4.5E8 pscbe2 = 1E-8 pvag = 0
+ delta = 0.01 fprout = 0 pdits = 1.4427E-15
+ pditsl = 0 pditsd = 0 lambda = 0
+ vtl = 0 lc = 0 xn = 0
+ alpha0 = 2.636988358999999E-5 walpha0 = 3.671447870068002E-11 alpha1 = 0
+ beta0 = 17.166379243999998 wbeta0 = 1.85538498868801E-6 aigbacc = 1
+ bigbacc = 0 cigbacc = 0 nigbacc = 1
+ aigbinv = 0.35 bigbinv = 0.03 cigbinv = 6E-3
+ eigbinv = 1.1 nigbinv = 3 aigc = 0.43
+ bigc = 0.054 cigc = 0.075 aigsd = 0.43
+ bigsd = 0.054 cigsd = 0.075 dlcig = 0
+ nigc = 1 poxedge = 1 pigcd = 1
+ ntox = 1 toxref = 4.148E-9 agidl = 0
+ bgidl = 2.3E9 cgidl = 0.5 egidl = 0.8
+ noia = 9E41 noib = 1E27 noic = 8E11
+ em = 4.1E7 af = 1 ef = 1.2
+ kf = 0 lintnoi = -3E-7 tnoia = 2.5E7
+ tnoib = 9.9E6 ntnoi = 1 rnoia = 0.912
+ rnoib = 0.26 xpart = 0 cgso = {2.392894381E-10/sw_func_tox_lv_ratio}
+ cgdo = {2.392894381E-10/sw_func_tox_lv_ratio} cgbo = {1E-14/sw_func_tox_lv_ratio} ckappas = 0.6
+ cf = 1E-14 clc = 1E-7 cle = 0.6
+ dlc = 1.21071E-8 dwc = 2.6E-8 vfbcv = -1
+ noff = 3.8661 voffcv = -0.16994 acde = 0.38008
+ moin = 23.81 cgsl = {2.310725E-11/sw_func_tox_lv_ratio} cgdl = {2.310725E-11/sw_func_tox_lv_ratio}
+ ijthsrev = 0.1 ijthsfwd = 0.1 xjbvs = 1
+ bvs = 11.9 jss = 2.75E-3 jsws = 6E-10
+ cjs = {1.210E-03*sw_func_nsd_pw_cj} mjs = 0.42197 mjsws = 1E-3
+ cjsws = {3.230311424E-11*sw_func_nsd_pw_cj} cjswgs = {1.795291232E-10*sw_func_nsd_pw_cj} mjswgs = 0.8
+ pbs = 0.7477 pbsws = 0.1 pbswgs = 0.79644
+ xrcrg1 = 12 xrcrg2 = 1 rbpb = 50
+ rbpd = 50 rbps = 50 rbdb = 50
+ rbsb = 50 gbmin = 1E-12 tnom = 30
+ ute = -1.1024166 wute = -4.675038631999987E-7 kt1 = -0.25142102
+ wkt1 = -1.290923304000036E-8 kt1l = 0 kt2 = -0.03455734
+ wkt2 = -6.564016799999985E-10 ua1 = 4.164049599999999E-9 wua1 = -6.129333020799997E-15
+ ub1 = -5.018905599999999E-18 wub1 = 8.638246108799998E-24 uc1 = 2.272055999999987E-12
+ wuc1 = -1.44729277088E-16 at = -3.009724899999999E5 wat = 1.82614594052
+ prt = 0 njs = 1.2928 xtis = 2
+ tpb = 1.2287E-3 tpbsw = 0 tpbswg = 0
+ tcj = 7.92E-4 tcjsw = 1E-5 tcjswg = 0
+ tvoff = 0 tvfbsdoff = 0 saref = 3E-6
+ sbref = 3E-6 wlod = 0 ku0 = -2.7E-8
+ kvsat = 0.2 kvth0 = 7.9E-9 tku0 = 0
+ llodku0 = 0 wlodku0 = 1 llodvth = 0
+ wlodvth = 1 lku0 = 0 wku0 = 0
+ pku0 = 0 lkvth0 = 0 wkvth0 = 3E-7
+ pkvth0 = 0 stk2 = 0 lodk2 = 1
+ steta0 = 0 lodeta0 = 1

.model nlowvt_model.18 nmos
+ level = 54 lmin = 4E-6 lmax = 8E-6 wmin = 3E-6
+ wmax = 5E-6 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 4.148E-9
+ toxm = 4.148E-9 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 9.999999999999999E22 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {2.6E-8+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {1.2025E-8-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = -1.33E-8 dwb = -1.08E-8 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = 0.428625 vfb = 0
+ k1 = 0.24736776 wk1 = 7.567582035200001E-7 k2 = 0.05125898698
+ wk2 = -2.958932598450399E-7 k3 = 1.65 k3b = 1.6
+ w0 = 1E-7 lpe0 = 2.3802E-7 lpeb = -4.9152E-8
+ vbm = -3 dvtp0 = 0 dvtp1 = 0
+ dvt0 = 0.07665 dvt1 = 0.1252 dvt2 = -0.05637
+ dvt0w = 0 dvt1w = 5.3E6 dvt2w = -0.032
+ vfbsdoff = 0 u0 = 0.0320233044 wu0 = 1.855428748799963E-9
+ ua = -1.508486209E-9 wua = 1.201240601131999E-15 ub = 2.94084734E-18
+ wub = -1.385080478320001E-24 uc = 7.254987096200001E-11 wuc = -1.043469351997604E-17
+ ud = 0 up = 0 lp = 1
+ eu = 1.67 vsat = 3.5078784E5 wvsat = -0.53358163232
+ a0 = 2.2794517696 wa0 = -1.754929275580798E-6 ags = 0.565636564
+ wags = -8.960612267200013E-8 b0 = 0 b1 = 0
+ keta = 0 a1 = 0 a2 = 0.38689047
+ rdsw = 103.65 rdswmin = 0 rdw = 0
+ rdwmin = 0 rsw = 0 rswmin = 0
+ prwb = 0 prwg = 0 wr = 1
+ voff = -0.1249454834 wvoff = 2.989617918319996E-8 voffl = 0
+ minv = 0 nfactor = 0.5601947258 wnfactor = 2.282660910261599E-6
+ eta0 = 0.08 etab = -0.07 dsub = 0.56
+ cit = 1.737E-5 wcit = -3.646676E-11 cdsc = 3.8556E-37
+ cdscb = -1.1484E-4 cdscd = 4.7984E-6 pclm = -0.125464596
+ wpclm = 9.59469629008E-7 pdiblc1 = 0.39 pdiblc2 = 6.403487E-3
+ wpdiblc2 = 9.08022323999997E-10 pdiblcb = 0 drout = 3.4946
+ pscbe1 = 4.5E8 pscbe2 = 1E-8 pvag = 0
+ delta = 0.01 fprout = 0 pdits = 1.4427E-15
+ pditsl = 0 pditsd = 0 lambda = 0
+ vtl = 0 lc = 0 xn = 0
+ alpha0 = 2.636988358999999E-5 walpha0 = 3.671447870068002E-11 alpha1 = 0
+ beta0 = 17.166379243999998 wbeta0 = 1.85538498868801E-6 aigbacc = 1
+ bigbacc = 0 cigbacc = 0 nigbacc = 1
+ aigbinv = 0.35 bigbinv = 0.03 cigbinv = 6E-3
+ eigbinv = 1.1 nigbinv = 3 aigc = 0.43
+ bigc = 0.054 cigc = 0.075 aigsd = 0.43
+ bigsd = 0.054 cigsd = 0.075 dlcig = 0
+ nigc = 1 poxedge = 1 pigcd = 1
+ ntox = 1 toxref = 4.148E-9 agidl = 0
+ bgidl = 2.3E9 cgidl = 0.5 egidl = 0.8
+ noia = 9E41 noib = 1E27 noic = 8E11
+ em = 4.1E7 af = 1 ef = 1.2
+ kf = 0 lintnoi = -3E-7 tnoia = 2.5E7
+ tnoib = 9.9E6 ntnoi = 1 rnoia = 0.912
+ rnoib = 0.26 xpart = 0 cgso = {2.392894381E-10/sw_func_tox_lv_ratio}
+ cgdo = {2.392894381E-10/sw_func_tox_lv_ratio} cgbo = {1E-14/sw_func_tox_lv_ratio} ckappas = 0.6
+ cf = 1E-14 clc = 1E-7 cle = 0.6
+ dlc = 1.21071E-8 dwc = 2.6E-8 vfbcv = -1
+ noff = 3.8661 voffcv = -0.16994 acde = 0.38008
+ moin = 23.81 cgsl = {2.310725E-11/sw_func_tox_lv_ratio} cgdl = {2.310725E-11/sw_func_tox_lv_ratio}
+ ijthsrev = 0.1 ijthsfwd = 0.1 xjbvs = 1
+ bvs = 11.9 jss = 2.75E-3 jsws = 6E-10
+ cjs = {1.210E-03*sw_func_nsd_pw_cj} mjs = 0.42197 mjsws = 1E-3
+ cjsws = {3.230311424E-11*sw_func_nsd_pw_cj} cjswgs = {1.795291232E-10*sw_func_nsd_pw_cj} mjswgs = 0.8
+ pbs = 0.7477 pbsws = 0.1 pbswgs = 0.79644
+ xrcrg1 = 12 xrcrg2 = 1 rbpb = 50
+ rbpd = 50 rbps = 50 rbdb = 50
+ rbsb = 50 gbmin = 1E-12 tnom = 30
+ ute = -1.1024166 wute = -4.675038631999987E-7 kt1 = -0.25142102
+ wkt1 = -1.290923304000036E-8 kt1l = 0 kt2 = -0.03455734
+ wkt2 = -6.564016799999985E-10 ua1 = 4.164049599999999E-9 wua1 = -6.129333020799997E-15
+ ub1 = -5.018905599999999E-18 wub1 = 8.638246108799998E-24 uc1 = 2.272055999999987E-12
+ wuc1 = -1.44729277088E-16 at = -3.009724899999999E5 wat = 1.82614594052
+ prt = 0 njs = 1.2928 xtis = 2
+ tpb = 1.2287E-3 tpbsw = 0 tpbswg = 0
+ tcj = 7.92E-4 tcjsw = 1E-5 tcjswg = 0
+ tvoff = 0 tvfbsdoff = 0 saref = 3E-6
+ sbref = 3E-6 wlod = 0 ku0 = -2.7E-8
+ kvsat = 0.2 kvth0 = 7.9E-9 tku0 = 0
+ llodku0 = 0 wlodku0 = 1 llodvth = 0
+ wlodvth = 1 lku0 = 0 wku0 = 0
+ pku0 = 0 lkvth0 = 0 wkvth0 = 3E-7
+ pkvth0 = 0 stk2 = 0 lodk2 = 1
+ steta0 = 0 lodeta0 = 1

.model nlowvt_model.19 nmos
+ level = 54 lmin = 2E-6 lmax = 4E-6 wmin = 3E-6
+ wmax = 5E-6 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 4.148E-9
+ toxm = 4.148E-9 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 9.999999999999999E22 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {2.6E-8+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {1.2025E-8-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = -1.33E-8 dwb = -1.08E-8 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = 0.442642682944778 lvth0 = -5.668971433344858E-8
+ wvth0 = -6.112888885114476E-8 pvth0 = 2.458640115080716E-13 vfb = 0
+ k1 = -0.0744791057355 lk1 = 1.279647045821062E-6 wk1 = 1.884946736685255E-6
+ pk1 = -4.485621198438394E-12 k2 = 0.17482886896565 lk2 = -4.913076722808472E-7
+ wk2 = -7.427456293140361E-7 pk2 = 1.776662678390255E-12 k3 = 1.65
+ k3b = 1.6 w0 = 1E-7 lpe0 = 2.3802E-7
+ lpeb = -4.9152E-8 vbm = -3 dvtp0 = 0
+ dvtp1 = 0 dvt0 = 0.07665 dvt1 = 0.1252
+ dvt2 = -0.05637 dvt0w = 0 dvt1w = 5.3E6
+ dvt2w = -0.032 vfbsdoff = 0 u0 = 0.030324367217109
+ lu0 = 6.754889292315424E-9 wu0 = 8.095088826778602E-9 pu0 = -2.480857648703916E-14
+ ua = -1.738562671546166E-9 lua = 9.1477251126043E-16 wua = 2.271143428580736E-15
+ pua = -4.253880146794802E-21 ub = 3.177572216166501E-18 lub = -9.412062713941993E-25
+ wub = -2.473926165530846E-24 pub = 4.32919601006596E-30 uc = 3.828139193978195E-11
+ luc = 1.362497591683878E-16 wuc = 3.26211299185588E-17 puc = -1.711878012004426E-22
+ ud = 0 up = 0 lp = 1
+ eu = 1.67 vsat = 6.3403080572355E5 lvsat = -1.126159869568549
+ wvsat = -0.985066009419925 pvsat = 1.795079309130449E-6 a0 = 2.521388656899489
+ la0 = -9.61928967058407E-7 wa0 = -2.930506482867625E-6 pa0 = 4.674036197312057E-12
+ ags = 0.287638040281599 lags = 1.105308230378174E-6 wags = -2.882112330099957E-6
+ pags = 1.110286505542318E-11 b0 = 0 b1 = 0
+ keta = 0.1612533868785 lketa = -6.411354035595723E-7 wketa = 2.58034306525182E-7
+ pketa = -1.025931501028797E-12 a1 = 0 a2 = 0.38689047
+ rdsw = 103.65 rdswmin = 0 rdw = 0
+ rdwmin = 0 rsw = 0 rswmin = 0
+ prwb = 0 prwg = 0 wr = 1
+ voff = -0.147918757298952 lvoff = 9.134058835854014E-8 wvoff = 1.066460733693769E-7
+ pvoff = -3.051537417895301E-13 voffl = 0 minv = 0
+ nfactor = -0.74262359224006 lnfactor = 5.179940491611377E-6 wnfactor = 6.182181129403963E-6
+ pnfactor = -1.550429741529908E-11 eta0 = 0.1585440125 leta0 = -3.122870664993751E-7
+ etab = -0.138652859865576 letab = 2.72960338182535E-7 wetab = -5.642023513242845E-11
+ petab = 2.243240338747788E-16 dsub = 0.584658173221702 ldsub = -9.803966382082431E-8
+ wdsub = 5.557500524720652E-7 pdsub = -2.209634421126307E-12 cit = 2.959125075000001E-5
+ lcit = -4.859108191946251E-11 wcit = -7.249500721100002E-11 pcit = 1.432465094985755E-16
+ cdsc = 3.8556E-37 cdscb = -1.1484E-4 cdscd = 4.7984E-6
+ pclm = -0.102331556565 lpclm = -9.197580814158841E-8 wpclm = 9.385732456256198E-7
+ ppclm = 8.308297550917417E-14 pdiblc1 = 0.39 pdiblc2 = 2.88673545128E-3
+ lpdiblc2 = 1.398242832013329E-8 wpdiblc2 = 7.571806928146559E-9 ppdiblc2 = -2.649487439685652E-14
+ pdiblcb = 0 drout = 3.4946 pscbe1 = 4.5E8
+ pscbe2 = 1E-8 pvag = 0 delta = 0.01
+ fprout = 0 pdits = 1.4427E-15 pditsl = 0
+ pditsd = 0 lambda = 0 vtl = 0
+ lc = 0 xn = 0 alpha0 = -5.63177008121598E-5
+ lalpha0 = 3.287617012037672E-10 walpha0 = -2.006196771192116E-11 palpha0 = 2.257403121141816E-16
+ alpha1 = 0 beta0 = 13.286509806054195 lbeta0 = 1.542616689180062E-5
+ wbeta0 = 2.593762298329145E-6 pbeta0 = -2.935751264267672E-12 aigbacc = 1
+ bigbacc = 0 cigbacc = 0 nigbacc = 1
+ aigbinv = 0.35 bigbinv = 0.03 cigbinv = 6E-3
+ eigbinv = 1.1 nigbinv = 3 aigc = 0.43
+ bigc = 0.054 cigc = 0.075 aigsd = 0.43
+ bigsd = 0.054 cigsd = 0.075 dlcig = 0
+ nigc = 1 poxedge = 1 pigcd = 1
+ ntox = 1 toxref = 4.148E-9 agidl = 0
+ bgidl = 2.3E9 cgidl = 0.5 egidl = 0.8
+ noia = 9E41 noib = 1E27 noic = 8E11
+ em = 4.1E7 af = 1 ef = 1.2
+ kf = 0 lintnoi = -3E-7 tnoia = 2.5E7
+ tnoib = 9.9E6 ntnoi = 1 rnoia = 0.912
+ rnoib = 0.26 xpart = 0 cgso = {2.392894381E-10/sw_func_tox_lv_ratio}
+ cgdo = {2.392894381E-10/sw_func_tox_lv_ratio} cgbo = {1E-14/sw_func_tox_lv_ratio} ckappas = 0.6
+ cf = 1E-14 clc = 1E-7 cle = 0.6
+ dlc = 1.21071E-8 dwc = 2.6E-8 vfbcv = -1
+ noff = 3.8661 voffcv = -0.16994 acde = 0.38008
+ moin = 23.81 cgsl = {2.310725E-11/sw_func_tox_lv_ratio} cgdl = {2.310725E-11/sw_func_tox_lv_ratio}
+ ijthsrev = 0.1 ijthsfwd = 0.1 xjbvs = 1
+ bvs = 11.9 jss = 2.75E-3 jsws = 6E-10
+ cjs = {1.210E-03*sw_func_nsd_pw_cj} mjs = 0.42197 mjsws = 1E-3
+ cjsws = {3.230311424E-11*sw_func_nsd_pw_cj} cjswgs = {1.795291232E-10*sw_func_nsd_pw_cj} mjswgs = 0.8
+ pbs = 0.7477 pbsws = 0.1 pbswgs = 0.79644
+ xrcrg1 = 12 xrcrg2 = 1 rbpb = 50
+ rbpd = 50 rbps = 50 rbdb = 50
+ rbsb = 50 gbmin = 1E-12 tnom = 30
+ ute = -0.93936831942 lute = -6.482718111720506E-7 wute = -1.095836494559838E-6
+ pute = 2.498219125655155E-12 kt1 = -0.2221776120635 lkt1 = -1.162703277851275E-7
+ wkt1 = -1.059341673388026E-7 pkt1 = 3.698624875253228E-13 kt1l = 0
+ kt2 = -0.0680812997962 lkt2 = 1.332895879517014E-7 wkt2 = 1.024420305389976E-7
+ pkt2 = -4.099142115811236E-13 ua1 = 5.096081108409998E-9 lua1 = -3.705710675862736E-15
+ wua1 = -9.295495385702674E-15 pua1 = 1.25885032547348E-20 ub1 = -6.58926854629E-18
+ lub1 = 6.243684556301727E-24 wub1 = 1.446473424776292E-23 pub1 = -2.316582551610963E-29
+ uc1 = 2.317189452855E-11 luc1 = -8.309671299758839E-17 wuc1 = -1.869327658709654E-16
+ puc1 = 1.677989612266313E-22 at = -6.784322037082E5 lat = 1.500760948718118
+ wat = 3.742041659407674 pat = -7.617505583511448E-6 prt = 0
+ njs = 1.2928 xtis = 2 tpb = 1.2287E-3
+ tpbsw = 0 tpbswg = 0 tcj = 7.92E-4
+ tcjsw = 1E-5 tcjswg = 0 tvoff = 0
+ tvfbsdoff = 0 saref = 3E-6 sbref = 3E-6
+ wlod = 0 ku0 = -2.7E-8 kvsat = 0.2
+ kvth0 = 7.9E-9 tku0 = 0 llodku0 = 0
+ wlodku0 = 1 llodvth = 0 wlodvth = 1
+ lku0 = 0 wku0 = 0 pku0 = 0
+ lkvth0 = 0 wkvth0 = 3E-7 pkvth0 = 0
+ stk2 = 0 lodk2 = 1 steta0 = 0
+ lodeta0 = 1

.model nlowvt_model.20 nmos
+ level = 54 lmin = 1E-6 lmax = 2E-6 wmin = 3E-6
+ wmax = 5E-6 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 4.148E-9
+ toxm = 4.148E-9 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 9.999999999999999E22 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {2.6E-8+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {1.2025E-8-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = -1.33E-8 dwb = -1.08E-8 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = 0.398811713900966 lvth0 = 2.991808894867145E-8
+ wvth0 = 1.027454623606307E-7 pvth0 = -7.79435127688362E-14 vfb = 0
+ k1 = 0.710430108482 lk1 = -2.71294316012008E-7 wk1 = -7.762219209489363E-7
+ pk1 = 7.727150106138865E-13 k2 = -0.12174872154293 lk2 = 9.471481768458248E-8
+ wk2 = 3.090287577896775E-7 pk2 = -3.015909218073283E-13 k3 = 1.65
+ k3b = 1.6 w0 = 1E-7 lpe0 = 2.3802E-7
+ lpeb = -4.9152E-8 vbm = -3 dvtp0 = 0
+ dvtp1 = 0 dvt0 = 0.07665 dvt1 = 0.1252
+ dvt2 = -0.05637 dvt0w = 0 dvt1w = 5.3E6
+ dvt2w = -0.032 vfbsdoff = 0 u0 = 0.036727439570295
+ lu0 = -5.897261523962404E-9 wu0 = -2.165706303893672E-9 pu0 = -4.533758348587284E-15
+ ua = -9.628326644889952E-10 lua = -6.180311961841872E-16 wua = -7.577906637394775E-17
+ pua = 3.835213571109048E-22 ub = 2.536206844822E-18 lub = 3.260996341139691E-25
+ wub = 8.900184657874563E-26 pub = -7.350215954619888E-31 uc = 1.337410924271E-10
+ luc = -5.237383600952822E-17 wuc = -8.787463824109068E-17 puc = 6.690581189461684E-23
+ ud = 0 up = 0 lp = 1
+ eu = 1.67 vsat = 6.041798509739997E4 lvsat = 7.270383347692483E-3
+ wvsat = -0.180936941487535 pvsat = 2.061604773494419E-7 a0 = 1.98243519102194
+ la0 = 1.030161338423378E-7 wa0 = 4.262030125333216E-7 pa0 = -1.958653930125444E-12
+ ags = -0.226038430210199 lags = 2.120307252246443E-6 wags = 5.050463432440066E-6
+ pags = -4.571508022567777E-12 b0 = 0 b1 = 0
+ keta = -0.180969781159 lketa = 3.508046532412607E-8 wketa = -3.997613609592677E-7
+ pketa = 2.738398481371014E-13 a1 = 0 a2 = 0.38689047
+ rdsw = 103.65 rdswmin = 0 rdw = 0
+ rdwmin = 0 rsw = 0 rswmin = 0
+ prwb = 0 prwg = 0 wr = 1
+ voff = -0.088953110847027 lvoff = -2.5172580748142E-8 wvoff = -9.053049606760238E-8
+ pvoff = 8.445730058946909E-14 voffl = 0 minv = 0
+ nfactor = 2.253322239797277 lnfactor = -7.398986752028012E-7 wnfactor = -4.318812439997797E-6
+ pnfactor = 5.245140828160332E-12 eta0 = 5.169974184659999E-4 leta0 = -3.358604901789242E-11
+ weta0 = 4.825967987623246E-11 peta0 = -9.535871445144154E-17 etab = -5.40780140278E-4
+ letab = 5.777424933331385E-11 wetab = 8.74293998875438E-11 petab = -5.991565244294003E-17
+ dsub = -0.227635633370691 ldsub = 1.507012283315414E-6 wdsub = 4.169434627720907E-7
+ pdsub = -1.935359540208643E-12 cit = 5E-6 cdsc = 3.8556E-37
+ cdscb = -1.1484E-4 cdscd = 4.7984E-6 pclm = -0.8247510153412
+ lpclm = 1.335488921427244E-6 wpclm = 3.242732341457857E-6 ppclm = -4.469820189900535E-12
+ pdiblc1 = 0.39 pdiblc2 = 9.676421495390001E-3 lpdiblc2 = 5.663481812741255E-10
+ wpdiblc2 = -2.008201670534972E-8 ppdiblc2 = 2.814769841175047E-14 pdiblcb = 0
+ drout = 3.4946 pscbe1 = 4.5E8 pscbe2 = 1E-8
+ pvag = 0 delta = 0.01 fprout = 0
+ pdits = 1.4427E-15 pditsl = 0 pditsd = 0
+ lambda = 0 vtl = 0 lc = 0
+ xn = 0 alpha0 = 1.410810632831775E-4 lalpha0 = -6.128838671041458E-11
+ walpha0 = 2.753271358239119E-10 palpha0 = -3.579337870174478E-16 alpha1 = 0
+ beta0 = 20.34658081183511 lbeta0 = 1.475819587927818E-6 wbeta0 = 5.20000728128849E-6
+ pbeta0 = -8.08556103834619E-12 aigbacc = 1 bigbacc = 0
+ cigbacc = 0 nigbacc = 1 aigbinv = 0.35
+ bigbinv = 0.03 cigbinv = 6E-3 eigbinv = 1.1
+ nigbinv = 3 aigc = 0.43 bigc = 0.054
+ cigc = 0.075 aigsd = 0.43 bigsd = 0.054
+ cigsd = 0.075 dlcig = 0 nigc = 1
+ poxedge = 1 pigcd = 1 ntox = 1
+ toxref = 4.148E-9 agidl = 0 bgidl = 2.3E9
+ cgidl = 0.5 egidl = 0.8 noia = 9E41
+ noib = 1E27 noic = 8E11 em = 4.1E7
+ af = 1 ef = 1.2 kf = 0
+ lintnoi = -3E-7 tnoia = 2.5E7 tnoib = 9.9E6
+ ntnoi = 1 rnoia = 0.912 rnoib = 0.26
+ xpart = 0 cgso = {2.392894381E-10/sw_func_tox_lv_ratio} cgdo = {2.392894381E-10/sw_func_tox_lv_ratio}
+ cgbo = {1E-14/sw_func_tox_lv_ratio} ckappas = 0.6 cf = 1E-14
+ clc = 1E-7 cle = 0.6 dlc = 1.21071E-8
+ dwc = 2.6E-8 vfbcv = -1 noff = 3.8661
+ voffcv = -0.16994 acde = 0.38008 moin = 23.81
+ cgsl = {2.310725E-11/sw_func_tox_lv_ratio} cgdl = {2.310725E-11/sw_func_tox_lv_ratio} ijthsrev = 0.1
+ ijthsfwd = 0.1 xjbvs = 1 bvs = 11.9
+ jss = 2.75E-3 jsws = 6E-10 cjs = {1.210E-03*sw_func_nsd_pw_cj}
+ mjs = 0.42197 mjsws = 1E-3 cjsws = {3.230311424E-11*sw_func_nsd_pw_cj}
+ cjswgs = {1.795291232E-10*sw_func_nsd_pw_cj} mjswgs = 0.8 pbs = 0.7477
+ pbsws = 0.1 pbswgs = 0.79644 xrcrg1 = 12
+ xrcrg2 = 1 rbpb = 50 rbpd = 50
+ rbps = 50 rbdb = 50 rbsb = 50
+ gbmin = 1E-12 tnom = 30 ute = -1.26415888698
+ lute = -6.501889201868656E-9 wute = -1.404424635829582E-7 pute = 6.10408290146388E-13
+ kt1 = -0.298329165073 lkt1 = 3.420133338399429E-8 wkt1 = 1.660226886732037E-7
+ pkt1 = -1.675106621116011E-13 kt1l = 0 kt2 = 0.054658237624
+ lkt2 = -1.092376010137428E-7 wkt2 = -3.11999577494352E-7 pkt2 = 4.090016838123736E-13
+ ua1 = 4.992482727259999E-9 lua1 = -3.501005454629396E-15 wua1 = -9.50304066256248E-15
+ pua1 = 1.299860234454593E-20 ub1 = -5.964041032829998E-18 lub1 = 5.008266251080435E-24
+ wub1 = 1.182405370078284E-23 pub1 = -1.794797278930432E-29 uc1 = -9.580199112109997E-11
+ luc1 = 1.519897363518375E-16 wuc1 = 2.235414222278026E-16 puc1 = -6.432775107471295E-22
+ at = 9.309106646429995E4 lat = -0.023730456979234 wat = -0.247462791180356
+ pat = 2.65555735627972E-7 prt = 0 njs = 1.2928
+ xtis = 2 tpb = 1.2287E-3 tpbsw = 0
+ tpbswg = 0 tcj = 7.92E-4 tcjsw = 1E-5
+ tcjswg = 0 tvoff = 0 tvfbsdoff = 0
+ saref = 3E-6 sbref = 3E-6 wlod = 0
+ ku0 = -2.7E-8 kvsat = 0.2 kvth0 = 7.9E-9
+ tku0 = 0 llodku0 = 0 wlodku0 = 1
+ llodvth = 0 wlodvth = 1 lku0 = 0
+ wku0 = 0 pku0 = 0 lkvth0 = 0
+ wkvth0 = 3E-7 pkvth0 = 0 stk2 = 0
+ lodk2 = 1 steta0 = 0 lodeta0 = 1

.model nlowvt_model.21 nmos
+ level = 54 lmin = 5E-7 lmax = 1E-6 wmin = 3E-6
+ wmax = 5E-6 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 4.148E-9
+ toxm = 4.148E-9 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 9.999999999999999E22 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {2.6E-8+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {1.2025E-8-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = -1.33E-8 dwb = -1.08E-8 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = 0.435585771958898 lvth0 = -5.97155301296763E-9
+ wvth0 = 2.767274848161202E-8 pvth0 = -4.676297658607877E-15 vfb = 0
+ k1 = 0.403113259874 lk1 = 2.863156238696971E-8 wk1 = 1.211309000634481E-7
+ pk1 = -1.0305647505315E-13 k2 = -7.948798447977806E-3 lk2 = -1.634821725993607E-8
+ wk2 = -4.202804133164503E-8 pk2 = 4.10229612951265E-14 k3 = 1.65
+ k3b = 1.6 w0 = 1E-7 lpe0 = 2.3802E-7
+ lpeb = -4.9152E-8 vbm = -3 dvtp0 = 0
+ dvtp1 = 0 dvt0 = 0.07665 dvt1 = 0.1252
+ dvt2 = -0.05637 dvt0w = 0 dvt1w = 5.3E6
+ dvt2w = -0.032 vfbsdoff = 0 u0 = 0.036967324866288
+ lu0 = -6.131377578586768E-9 wu0 = -2.542053285971301E-8 pu0 = 1.81617896285646E-14
+ ua = -1.067094938118585E-9 lua = -5.162764302353894E-16 wua = -1.890204264228053E-15
+ pua = 2.154309628956619E-21 ub = 2.603257519366E-18 lub = 2.606615282927521E-25
+ wub = 1.379682238197034E-24 pub = -1.994661123661857E-30 uc = 9.266922486547523E-11
+ luc = -1.228974686276054E-17 wuc = 1.4172176093379E-17 puc = -3.268677655510885E-23
+ ud = 0 up = 0 lp = 1
+ eu = 1.67 vsat = -7.229307141947998E4 lvsat = 0.136789738955342
+ wvsat = 0.188356394960147 pvsat = -1.542513543566736E-7 a0 = 2.9242970018204
+ la0 = -8.16193900406419E-7 wa0 = -4.760637528898537E-6 pa0 = 3.103443096284979E-12
+ ags = 4.810877487260999 lags = -2.795470837409572E-6 wags = -4.534681912709828E-6
+ pags = 4.783114577031262E-12 b0 = 0 b1 = 0
+ keta = -0.300055605122154 lketa = 1.513022752209666E-7 wketa = -1.4858944878758E-7
+ pketa = 2.870862045314276E-14 a1 = 0 a2 = 0.38689047
+ rdsw = 103.65 rdswmin = 0 rdw = 0
+ rdwmin = 0 rsw = 0 rswmin = 0
+ prwb = 0 prwg = 0 wr = 1
+ voff = -0.11028928224414 lvoff = -4.349544273129539E-9 wvoff = -3.105466535263914E-8
+ pvoff = 2.641186360320072E-14 voffl = 0 minv = 0
+ nfactor = 1.076563940394365 lnfactor = 4.085585870994718E-7 wnfactor = 5.152172091200447E-7
+ pnfactor = 5.273695921037745E-13 eta0 = 9.55986169068E-4 leta0 = -4.620171201679146E-10
+ weta0 = -1.659447774404643E-10 peta0 = 1.136941256667891E-16 etab = -9.308767654693791E-4
+ letab = 4.384890506888406E-10 wetab = 3.028407946484539E-10 petab = -2.701464031598507E-16
+ dsub = 1.617802573854576 ldsub = -2.940431350260853E-7 wdsub = -3.056887135432442E-6
+ pdsub = 1.45492543210907E-12 cit = 5E-6 cdsc = 3.8556E-37
+ cdscb = -1.1484E-4 cdscd = 4.7984E-6 pclm = 0.567970296698
+ lpclm = -2.373744305741311E-8 wpclm = -1.981712241597704E-6 ppclm = 6.289765009325392E-13
+ pdiblc1 = 0.39 pdiblc2 = 0.01204869069584 lpdiblc2 = -1.748867944905045E-9
+ wpdiblc2 = 9.964541003063691E-9 ppdiblc2 = -1.176239583775606E-15 pdiblcb = 0
+ drout = 3.4946 pscbe1 = 4.5E8 pscbe2 = 1E-8
+ pvag = 0 delta = 0.01 fprout = 0
+ pdits = 1.4427E-15 pditsl = 0 pditsd = 0
+ lambda = 0 vtl = 0 lc = 0
+ xn = 0 alpha0 = 2.488948285656302E-5 lalpha0 = 5.210878620693982E-11
+ walpha0 = -1.090653466631222E-10 palpha0 = 1.721405626577311E-17 alpha1 = 0
+ beta0 = 19.605310616645188 lbeta0 = 2.199262234923423E-6 wbeta0 = -4.672854344550807E-6
+ pbeta0 = 1.549858265391672E-12 aigbacc = 1 bigbacc = 0
+ cigbacc = 0 nigbacc = 1 aigbinv = 0.35
+ bigbinv = 0.03 cigbinv = 6E-3 eigbinv = 1.1
+ nigbinv = 3 aigc = 0.43 bigc = 0.054
+ cigc = 0.075 aigsd = 0.43 bigsd = 0.054
+ cigsd = 0.075 dlcig = 0 nigc = 1
+ poxedge = 1 pigcd = 1 ntox = 1
+ toxref = 4.148E-9 agidl = 0 bgidl = 2.3E9
+ cgidl = 0.5 egidl = 0.8 noia = 9E41
+ noib = 1E27 noic = 8E11 em = 4.1E7
+ af = 1 ef = 1.2 kf = 0
+ lintnoi = -3E-7 tnoia = 2.5E7 tnoib = 9.9E6
+ ntnoi = 1 rnoia = 0.912 rnoib = 0.26
+ xpart = 0 cgso = {2.392894381E-10/sw_func_tox_lv_ratio} cgdo = {2.392894381E-10/sw_func_tox_lv_ratio}
+ cgbo = {1E-14/sw_func_tox_lv_ratio} ckappas = 0.6 cf = 1E-14
+ clc = 1E-7 cle = 0.6 dlc = 1.21071E-8
+ dwc = 2.6E-8 vfbcv = -1 noff = 3.8661
+ voffcv = -0.16994 acde = 0.38008 moin = 23.81
+ cgsl = {2.310725E-11/sw_func_tox_lv_ratio} cgdl = {2.310725E-11/sw_func_tox_lv_ratio} ijthsrev = 0.1
+ ijthsfwd = 0.1 xjbvs = 1 bvs = 11.9
+ jss = 2.75E-3 jsws = 6E-10 cjs = {1.210E-03*sw_func_nsd_pw_cj}
+ mjs = 0.42197 mjsws = 1E-3 cjsws = {3.230311424E-11*sw_func_nsd_pw_cj}
+ cjswgs = {1.795291232E-10*sw_func_nsd_pw_cj} mjswgs = 0.8 pbs = 0.7477
+ pbsws = 0.1 pbswgs = 0.79644 xrcrg1 = 12
+ xrcrg2 = 1 rbpb = 50 rbpd = 50
+ rbps = 50 rbdb = 50 rbsb = 50
+ gbmin = 1E-12 tnom = 30 ute = -2.18448393852
+ lute = 8.916893448485938E-7 wute = 4.401989973956959E-6 pute = -3.822778647270694E-12
+ kt1 = -0.25104520423 lkt1 = -1.194544820073154E-8 wkt1 = -6.080908810196002E-8
+ pkt1 = 5.386581043211993E-14 kt1l = 0 kt2 = -0.0656849655074
+ lkt2 = 8.211348082347034E-9 wkt2 = 1.430364178846152E-7 pkt2 = -3.509069587772941E-14
+ ua1 = -2.505674732577999E-9 lua1 = 3.816821318299498E-15 wua1 = 2.209302550319594E-14
+ pua1 = -1.7837578429926E-20 ub1 = 4.297623203039997E-18 lub1 = -5.006604959916886E-24
+ wub1 = -3.009031333500191E-23 pub1 = 2.29583537192698E-29 uc1 = 1.783454618679999E-10
+ luc1 = -1.155644703928745E-16 wuc1 = -1.031119387775664E-15 puc1 = 5.812087067757535E-22
+ at = 1.166976457308E5 lat = -0.046769298014374 wat = -0.101842282887998
+ pat = 1.234374005600452E-7 prt = 0 njs = 1.2928
+ xtis = 2 tpb = 1.2287E-3 tpbsw = 0
+ tpbswg = 0 tcj = 7.92E-4 tcjsw = 1E-5
+ tcjswg = 0 tvoff = 0 tvfbsdoff = 0
+ saref = 2.74E-6 sbref = 2.74E-6 wlod = 0
+ ku0 = -2.7E-8 kvsat = 0.2 kvth0 = 7.9E-9
+ tku0 = 0 llodku0 = 0 wlodku0 = 1
+ llodvth = 0 wlodvth = 1 lku0 = 0
+ wku0 = 0 pku0 = 0 lkvth0 = 0
+ wkvth0 = 3E-7 pkvth0 = 0 stk2 = 0
+ lodk2 = 1 steta0 = 0 lodeta0 = 1

.model nlowvt_model.22 nmos
+ level = 54 lmin = 2.5E-7 lmax = 5E-7 wmin = 3E-6
+ wmax = 5E-6 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 4.148E-9
+ toxm = 4.148E-9 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 9.999999999999999E22 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {2.6E-8+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {1.2025E-8-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = -1.33E-8 dwb = -1.08E-8 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = 0.496857864570564 lvth0 = -3.513400549148992E-8
+ wvth0 = -3.446829301070315E-9 pvth0 = 1.013506538705978E-14 vfb = 0
+ k1 = 0.323905458464248 lk1 = 6.63305154679412E-8 wk1 = -1.089993458570988E-7
+ pk1 = 6.474015492734238E-15 k2 = -7.108015765796118E-4 lk2 = -1.979314187087803E-8
+ wk2 = 5.095966737545354E-8 pk2 = -3.234538664017061E-15 k3 = 1.65
+ k3b = 1.6 w0 = 1E-7 lpe0 = 2.3802E-7
+ lpeb = -4.9152E-8 vbm = -3 dvtp0 = 0
+ dvtp1 = 0 dvt0 = 0.07665 dvt1 = 0.1252
+ dvt2 = -0.05637 dvt0w = 0 dvt1w = 5.3E6
+ dvt2w = -0.032 vfbsdoff = 0 u0 = 0.017364276374536
+ lu0 = 3.198693351062777E-9 wu0 = 5.428873055127782E-8 pu0 = -1.977583429189648E-14
+ ua = -3.082184600420022E-9 lua = 4.428054945369799E-16 wua = 7.558705165754755E-15
+ pua = -2.342898814243698E-21 ub = 4.066423803696958E-18 lub = -4.357324647345676E-25
+ wub = -6.952680892228552E-24 pub = 1.9711271082642E-30 uc = 5.184868431814318E-11
+ luc = 7.138789410742147E-18 wuc = -8.011843347974104E-18 puc = -2.212829250199687E-23
+ ud = 0 up = 0 lp = 1
+ eu = 1.67 vsat = 2.72847170687976E5 lvsat = -0.027479759275702
+ wvsat = -0.288069899400905 pvsat = 7.250374044446934E-8 a0 = 1.05959741226524
+ la0 = 7.130986924235895E-8 wa0 = 3.032500689231592E-6 pa0 = -6.057010386340563E-13
+ ags = -2.022934789390799 lags = 4.57082115662851E-7 wags = 1.049933088270808E-5
+ pags = -2.37232381294789E-12 b0 = 0 b1 = 0
+ keta = 0.068806221124116 lketa = -2.4257510980946E-8 wketa = -1.822168822330823E-7
+ pketa = 4.471359740152955E-14 a1 = 0 a2 = 0.38689047
+ rdsw = 103.65 rdswmin = 0 rdw = 0
+ rdwmin = 0 rsw = 0 rswmin = 0
+ prwb = 0 prwg = 0 wr = 1
+ voff = -0.124751659736996 lvoff = 2.533824294595249E-9 wvoff = 3.89785113251042E-8
+ pvoff = -6.92042683657122E-15 voffl = 0 minv = 0
+ nfactor = 1.407480749251519 lnfactor = 2.510587319239092E-7 wnfactor = 3.176531166779883E-6
+ pnfactor = -7.392827860444253E-13 eta0 = 2.888320834652441E-3 leta0 = -1.381711804252828E-9
+ weta0 = -3.032446535115684E-8 peta0 = 1.446764199272709E-14 etab = 0.100956404709422
+ letab = -4.805476256728549E-8 wetab = -2.485946575733537E-7 petab = 1.181926179450908E-13
+ dsub = 1.496608150182892 ldsub = -2.363606490795475E-7 wdsub = 4.965392506544023E-7
+ pdsub = -2.363278563489627E-13 cit = 5E-6 cdsc = 3.8556E-37
+ cdscb = -1.1484E-4 cdscd = 4.7984E-6 pclm = 0.591445922776808
+ lpclm = -3.491066728962175E-8 wpclm = -1.058053604643646E-6 ppclm = 1.893611726742552E-13
+ pdiblc1 = 0.39 pdiblc2 = 5.367275584320002E-3 lpdiblc2 = 1.431151577422895E-9
+ wpdiblc2 = -1.110316569753716E-10 ppdiblc2 = 3.619229223769985E-15 pdiblcb = 0
+ drout = 3.4946 pscbe1 = 4.5E8 pscbe2 = 1E-8
+ pvag = 0 delta = 0.01 fprout = 0
+ pdits = 1.4427E-15 pditsl = 0 pditsd = 0
+ lambda = 0 vtl = 0 lc = 0
+ xn = 0 alpha0 = -1.189520411187396E-3 lalpha0 = 6.30107175277162E-10
+ walpha0 = -1.232694073215109E-9 palpha0 = 5.52005148668191E-16 alpha1 = 0
+ beta0 = 18.522351424777604 lbeta0 = 2.714696662292801E-6 wbeta0 = -2.518302275134774E-6
+ pbeta0 = 5.243992079531106E-13 aigbacc = 1 bigbacc = 0
+ cigbacc = 0 nigbacc = 1 aigbinv = 0.35
+ bigbinv = 0.03 cigbinv = 6E-3 eigbinv = 1.1
+ nigbinv = 3 aigc = 0.43 bigc = 0.054
+ cigc = 0.075 aigsd = 0.43 bigsd = 0.054
+ cigsd = 0.075 dlcig = 0 nigc = 1
+ poxedge = 1 pigcd = 1 ntox = 1
+ toxref = 4.148E-9 agidl = 0 bgidl = 2.3E9
+ cgidl = 0.5 egidl = 0.8 noia = 9E41
+ noib = 1E27 noic = 8E11 em = 4.1E7
+ af = 1 ef = 1.2 kf = 0
+ lintnoi = -3E-7 tnoia = 2.5E7 tnoib = 9.9E6
+ ntnoi = 1 rnoia = 0.912 rnoib = 0.26
+ xpart = 0 cgso = {2.392894381E-10/sw_func_tox_lv_ratio} cgdo = {2.392894381E-10/sw_func_tox_lv_ratio}
+ cgbo = {1E-14/sw_func_tox_lv_ratio} ckappas = 0.6 cf = 1E-14
+ clc = 1E-7 cle = 0.6 dlc = 1.21071E-8
+ dwc = 2.6E-8 vfbcv = -1 noff = 3.8661
+ voffcv = -0.16994 acde = 0.38008 moin = 23.81
+ cgsl = {2.310725E-11/sw_func_tox_lv_ratio} cgdl = {2.310725E-11/sw_func_tox_lv_ratio} ijthsrev = 0.1
+ ijthsfwd = 0.1 xjbvs = 1 bvs = 11.9
+ jss = 2.75E-3 jsws = 6E-10 cjs = {1.210E-03*sw_func_nsd_pw_cj}
+ mjs = 0.42197 mjsws = 1E-3 cjsws = {3.230311424E-11*sw_func_nsd_pw_cj}
+ cjswgs = {1.795291232E-10*sw_func_nsd_pw_cj} mjswgs = 0.8 pbs = 0.7477
+ pbsws = 0.1 pbswgs = 0.79644 xrcrg1 = 12
+ xrcrg2 = 1 rbpb = 50 rbpd = 50
+ rbps = 50 rbdb = 50 rbsb = 50
+ gbmin = 1E-12 tnom = 30 ute = -0.968759065472
+ lute = 3.130650915213983E-7 wute = -1.292736956428544E-6 pute = -1.112373364753714E-12
+ kt1 = -0.337465445036 lkt1 = 2.91862654108842E-8 wkt1 = 2.667952942781282E-7
+ pkt1 = -1.02057495361683E-13 kt1l = 0 kt2 = -0.0589458429632
+ lkt2 = 5.003862707435037E-9 wkt2 = 8.338866262031357E-8 pkt2 = -6.701346759685052E-15
+ ua1 = 4.841665203606001E-9 lua1 = 3.198548756727237E-16 wua1 = -1.265257574568249E-14
+ pua1 = -1.30040951552231E-21 ub1 = -6.468168265179201E-18 lub1 = 1.173734893820403E-25
+ wub1 = 1.853099252754668E-23 pub1 = -1.829568060102033E-31 uc1 = -1.628909896484E-10
+ luc1 = 4.684701870635596E-17 wuc1 = 5.605370342458832E-16 puc1 = -1.763401672854017E-22
+ at = 1.415265163200002E3 lat = 8.099351016774956E-3 wat = 0.248894995829286
+ pat = -4.349600724544645E-8 prt = 0 njs = 1.2928
+ xtis = 2 tpb = 1.2287E-3 tpbsw = 0
+ tpbswg = 0 tcj = 7.92E-4 tcjsw = 1E-5
+ tcjswg = 0 tvoff = 0 tvfbsdoff = 0
+ saref = 1.74E-6 sbref = 1.74E-6 wlod = 0
+ ku0 = -2.7E-8 kvsat = 0.2 kvth0 = 7.9E-9
+ tku0 = 0 llodku0 = 0 wlodku0 = 1
+ llodvth = 0 wlodvth = 1 lku0 = 0
+ wku0 = 0 pku0 = 0 lkvth0 = 0
+ wkvth0 = 3E-7 pkvth0 = 0 stk2 = 0
+ lodk2 = 1 steta0 = 0 lodeta0 = 1

.model nlowvt_model.23 nmos
+ level = 54 lmin = 1.8E-7 lmax = 2.5E-7 wmin = 3E-6
+ wmax = 5E-6 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 4.148E-9
+ toxm = 4.148E-9 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 9.999999999999999E22 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {2.6E-8+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {1.2025E-8-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = -1.33E-8 dwb = -1.08E-8 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = 0.6285056731447 lvth0 = -6.487982783881587E-8
+ wvth0 = -1.778726033342598E-7 pvth0 = 4.954656902985895E-14 vfb = 0
+ k1 = 0.388689572027686 lk1 = 5.16925450082824E-8 wk1 = -7.703969145013177E-8
+ pk1 = -7.472684205199576E-16 k2 = -0.029712537587017 lk2 = -1.324019961931969E-8
+ wk2 = 4.646344384723484E-8 pk2 = -2.218616957816044E-15 k3 = 1.65
+ k3b = 1.6 w0 = 1E-7 lpe0 = 2.3802E-7
+ lpeb = -4.9152E-8 vbm = -3 dvtp0 = 0
+ dvtp1 = 0 dvt0 = 0.07665 dvt1 = 0.1252
+ dvt2 = -0.05637 dvt0w = 0 dvt1w = 5.3E6
+ dvt2w = -0.032 vfbsdoff = 0 u0 = 0.072401617509101
+ lu0 = -9.236993878292364E-9 wu0 = -1.280763908626624E-7 pu0 = 2.14295648915833E-14
+ ua = 2.37390778660094E-9 lua = -7.899985803104064E-16 wua = -1.199895433095317E-14
+ pua = 2.076154349037456E-21 ub = 7.773456225371493E-20 lub = 4.655118693695331E-25
+ wub = 8.405994915654333E-24 pub = -1.499165690526937E-30 uc = 2.004511687715672E-10
+ luc = -2.6437941951509E-17 wuc = -3.949819345649258E-16 puc = 6.530759960847336E-23
+ ud = 0 up = 0 lp = 1
+ eu = 1.67 vsat = 9.341722926778576E4 lvsat = 0.01306243598819
+ wvsat = 0.193639777927568 pvsat = -3.633856114789915E-8 a0 = 4.438941493481286
+ la0 = -6.922529259084065E-7 wa0 = 1.135607029968885E-6 pa0 = -1.770979163236476E-13
+ ags = -2.820889544571429 lags = 6.373799925959142E-7 wags = 8.189267359679998E-7
+ pags = -1.850364959919696E-13 b0 = 0 b1 = 0
+ keta = -0.023681121363479 lketa = -3.359995945873923E-9 wketa = 4.824522719017977E-7
+ pketa = -1.054683979752466E-13 a1 = 0 a2 = 0.38689047
+ rdsw = 103.65 rdswmin = 0 rdw = 0
+ rdwmin = 0 rsw = 0 rswmin = 0
+ prwb = 0 prwg = 0 wr = 1
+ voff = -0.172155676009154 lvoff = 1.324476177128939E-8 wvoff = 6.104012369754073E-8
+ pvoff = -1.190524815212326E-14 voffl = 0 minv = 0
+ nfactor = 1.12811809949543 lnfactor = 3.141807226362976E-7 wnfactor = 5.960916686820443E-7
+ pnfactor = -1.562324814492188E-13 eta0 = -0.248514655629256 leta0 = 5.542279072776725E-8
+ weta0 = 2.841310068693172E-7 peta0 = -5.658357195548901E-14 etab = -0.315616350797248
+ letab = 4.60698515394466E-8 wetab = 8.506424048765314E-7 petab = -1.301799963154607E-13
+ dsub = 0.8031454468433 ldsub = -7.96727512599666E-8 wdsub = -2.056927022236476E-6
+ pdsub = 3.406278480107312E-13 cit = 1.004254565381657E-5 lcit = -1.139363190479855E-12
+ wcit = -1.486542458745126E-11 pcit = 3.358842685534612E-18 cdsc = 3.8556E-37
+ cdscb = -1.1484E-4 cdscd = 4.7984E-6 pclm = 1.347875348282828
+ lpclm = -2.05825895982707E-7 wpclm = -1.913453618217721E-6 ppclm = 3.826388057413175E-13
+ pdiblc1 = -0.978741819110314 lpdiblc1 = 3.092672140279754E-7 wpdiblc1 = 4.825395803320558E-8
+ ppdiblc1 = -1.09029818176028E-14 pdiblc2 = 0.02233499984 lpdiblc2 = -2.402705718148E-9
+ wpdiblc2 = 1.59717948973943E-8 ppdiblc2 = -1.46854361898408E-17 pdiblcb = 0
+ drout = 3.4946 pscbe1 = 4.5E8 pscbe2 = 1E-8
+ pvag = 0 delta = 0.01 fprout = 0
+ pdits = 1.4427E-15 pditsl = 0 pditsd = 0
+ lambda = 0 vtl = 0 lc = 0
+ xn = 0 alpha0 = -1.179903264515041E-3 lalpha0 = 6.279341809865437E-10
+ walpha0 = 1.9024676636103E-8 palpha0 = -4.025147763102236E-15 alpha1 = 0
+ beta0 = 25.148567965537143 lbeta0 = 1.217503034908182E-6 wbeta0 = 2.76462006792908E-5
+ pbeta0 = -6.291270234599348E-12 aigbacc = 1 bigbacc = 0
+ cigbacc = 0 nigbacc = 1 aigbinv = 0.35
+ bigbinv = 0.03 cigbinv = 6E-3 eigbinv = 1.1
+ nigbinv = 3 aigc = 0.43 bigc = 0.054
+ cigc = 0.075 aigsd = 0.43 bigsd = 0.054
+ cigsd = 0.075 dlcig = 0 nigc = 1
+ poxedge = 1 pigcd = 1 ntox = 1
+ toxref = 4.148E-9 agidl = 0 bgidl = 2.3E9
+ cgidl = 0.5 egidl = 0.8 noia = 9E41
+ noib = 1E27 noic = 8E11 em = 4.1E7
+ af = 1 ef = 1.2 kf = 0
+ lintnoi = -3E-7 tnoia = 2.5E7 tnoib = 9.9E6
+ ntnoi = 1 rnoia = 0.912 rnoib = 0.26
+ xpart = 0 cgso = {2.392894381E-10/sw_func_tox_lv_ratio} cgdo = {2.392894381E-10/sw_func_tox_lv_ratio}
+ cgbo = {1E-14/sw_func_tox_lv_ratio} ckappas = 0.6 cf = 1E-14
+ clc = 1E-7 cle = 0.6 dlc = 1.21071E-8
+ dwc = 2.6E-8 vfbcv = -1 noff = 3.8661
+ voffcv = -0.16994 acde = 0.38008 moin = 23.81
+ cgsl = {2.310725E-11/sw_func_tox_lv_ratio} cgdl = {2.310725E-11/sw_func_tox_lv_ratio} ijthsrev = 0.1
+ ijthsfwd = 0.1 xjbvs = 1 bvs = 11.9
+ jss = 2.75E-3 jsws = 6E-10 cjs = {1.210E-03*sw_func_nsd_pw_cj}
+ mjs = 0.42197 mjsws = 1E-3 cjsws = {3.230311424E-11*sw_func_nsd_pw_cj}
+ cjswgs = {1.795291232E-10*sw_func_nsd_pw_cj} mjswgs = 0.8 pbs = 0.7477
+ pbsws = 0.1 pbswgs = 0.79644 xrcrg1 = 12
+ xrcrg2 = 1 rbpb = 50 rbpd = 50
+ rbps = 50 rbdb = 50 rbsb = 50
+ gbmin = 1E-12 tnom = 30 ute = 4.442520274828572
+ lute = -9.096134754195155E-7 wute = -1.787351423876606E-5 pute = 2.634053262190446E-12
+ kt1 = 0.037287405028571 lkt1 = -5.54891410612057E-8 wkt1 = -7.022401889385138E-7
+ pkt1 = 1.168960720711172E-13 kt1l = 0 kt2 = -0.018523558155714
+ lkt2 = -4.129552544816359E-9 wkt2 = 2.12817771259028E-8 pkt2 = 7.331704017777056E-15
+ ua1 = 1.852774133771857E-8 lua1 = -2.77251402683001E-15 wua1 = -5.433180081720292E-14
+ pua1 = 8.117011389387727E-21 ub1 = -1.750897826740286E-17 lub1 = 2.612044509384475E-24
+ wub1 = 5.069597246448076E-23 pub1 = -7.450634022760458E-30 uc1 = 1.238246698574286E-10
+ luc1 = -1.793638455898598E-17 wuc1 = -6.126844664545566E-16 puc1 = 8.874923079786265E-23
+ at = -1.060859756871428E5 lat = 0.03238925638691 wat = 0.386676399291411
+ pat = -7.462771535771359E-8 prt = 0 njs = 1.2928
+ xtis = 2 tpb = 1.2287E-3 tpbsw = 0
+ tpbswg = 0 tcj = 7.92E-4 tcjsw = 1E-5
+ tcjswg = 0 tvoff = 0 tvfbsdoff = 0
+ saref = 1.25E-6 sbref = 1.24E-6 wlod = 0
+ ku0 = -2.7E-8 kvsat = 0.2 kvth0 = 7.9E-9
+ tku0 = 0 llodku0 = 0 wlodku0 = 1
+ llodvth = 0 wlodvth = 1 lku0 = 0
+ wku0 = 0 pku0 = 0 lkvth0 = 0
+ wkvth0 = 3E-7 pkvth0 = 0 stk2 = 0
+ lodk2 = 1 steta0 = 0 lodeta0 = 1

.model nlowvt_model.24 nmos
+ level = 54 lmin = 1.5E-7 lmax = 1.8E-7 wmin = 3E-6
+ wmax = 5E-6 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 4.148E-9
+ toxm = 4.148E-9 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 9.999999999999999E22 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {2.6E-8+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {1.2025E-8-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = -1.33E-8 dwb = -1.08E-8 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = 0.099277746973334 lvth0 = 1.765326724760865E-8
+ wvth0 = 7.655841805092792E-7 pvth0 = -9.758551641054091E-14 vfb = 0
+ k1 = 0.649774817033333 lk1 = 1.09763010496517E-8 wk1 = 6.723372894524011E-7
+ pk1 = -1.1761260859227E-13 k2 = -0.098733935538344 lk2 = -2.476312608810332E-9
+ wk2 = -2.540592671771433E-7 pk2 = 4.464789982643572E-14 k3 = 1.65
+ k3b = 1.6 w0 = 1E-7 lpe0 = 2.3802E-7
+ lpeb = -4.9152E-8 vbm = -3 dvtp0 = 0
+ dvtp1 = 0 dvt0 = 0.07665 dvt1 = 0.1252
+ dvt2 = -0.05637 dvt0w = 0 dvt1w = 5.3E6
+ dvt2w = -0.032 vfbsdoff = 0 u0 = -0.011033820294267
+ lu0 = 3.774762647142885E-9 wu0 = 1.144781236558314E-7 pu0 = -1.639681164757581E-14
+ ua = -2.897502182198662E-9 lua = 3.207780432389142E-17 wua = 3.550265311192318E-15
+ pua = -3.487464541551317E-22 ub = 1.539304513773332E-18 lub = 2.375800354300488E-25
+ wub = 3.935677066516216E-24 pub = -8.020196219538478E-31 uc = 1.1844428752489E-10
+ luc = -1.36489688210897E-17 wuc = -9.571235145982243E-17 puc = 1.863650812323249E-23
+ ud = 0 up = 0 lp = 1
+ eu = 1.67 vsat = 2.536932152506E5 lvsat = -0.01193260402583
+ wvsat = -0.294654534331969 pvsat = 3.981093684897557E-8 a0 = 0
+ ags = 1.299373226666666 lags = -5.174986578666645E-9 wags = -1.776101390213335E-6
+ pags = 2.196581402860095E-13 b0 = 0 b1 = 0
+ keta = -0.27390493456858 lketa = 3.566240772346163E-8 wketa = 1.283985518736574E-6
+ pketa = -2.304675078191299E-13 a1 = 0 a2 = 0.38689047
+ rdsw = 103.65 rdswmin = 0 rdw = 0
+ rdwmin = 0 rsw = 0 rswmin = 0
+ prwb = 0 prwg = 0 wr = 1
+ voff = 0.192436447187606 lvoff = -4.361337984124543E-8 wvoff = -9.641714559517172E-7
+ pvoff = 1.479764976941785E-13 voffl = 0 minv = 0
+ nfactor = 4.845023331208994 lnfactor = -2.654706482494326E-7 wnfactor = -1.130307157837011E-5
+ pnfactor = 1.699442026928565E-12 eta0 = 0.408388617711613 leta0 = -4.70212747497413E-8
+ weta0 = -9.547189672136497E-7 peta0 = 1.366150815027496E-13 etab = 0.017989878941687
+ letab = -5.956039988340336E-9 wetab = -2.800355438539123E-7 petab = 4.614922978905194E-14
+ dsub = 0.427692705841534 ldsub = -2.112089630074114E-8 wdsub = 6.616692964317591E-7
+ pdsub = -8.333724788558005E-14 cit = 2.417577680776132E-5 lcit = -3.343440588937537E-12
+ wcit = -1.184136233626137E-10 pcit = 1.95071842845212E-17 cdsc = 3.8556E-37
+ cdscb = -1.1484E-4 cdscd = 4.7984E-6 pclm = -1.602861501766666
+ lpclm = 2.543415157825116E-7 wpclm = 5.8836283792748E-6 ppclm = -8.333161317676408E-13
+ pdiblc1 = 2.192949832828533 lpdiblc1 = -1.853580990918878E-7 wpdiblc1 = -3.562348816202517E-6
+ ppdiblc1 = 5.521705208244581E-13 pdiblc2 = 0.041682559433667 lpdiblc2 = -5.419957636780318E-9
+ wpdiblc2 = -6.373870604449342E-9 ppdiblc2 = 3.470121098822674E-15 pdiblcb = 0
+ drout = 3.4946 pscbe1 = 4.5E8 pscbe2 = 1E-8
+ pvag = 0 delta = 0.01 fprout = 0
+ pdits = 1.4427E-15 pditsl = 0 pditsd = 0
+ lambda = 0 vtl = 0 lc = 0
+ xn = 0 alpha0 = 0.010150693018288 lalpha0 = -1.139072309316621E-9
+ walpha0 = -2.571383118600234E-8 palpha0 = 2.951822531755092E-15 alpha1 = 0
+ beta0 = 41.390217479650005 lbeta0 = -1.315382206817717E-6 wbeta0 = -2.907290968156153E-5
+ pbeta0 = 2.554075026175573E-12 aigbacc = 1 bigbacc = 0
+ cigbacc = 0 nigbacc = 1 aigbinv = 0.35
+ bigbinv = 0.03 cigbinv = 6E-3 eigbinv = 1.1
+ nigbinv = 3 aigc = 0.43 bigc = 0.054
+ cigc = 0.075 aigsd = 0.43 bigsd = 0.054
+ cigsd = 0.075 dlcig = 0 nigc = 1
+ poxedge = 1 pigcd = 1 ntox = 1
+ toxref = 4.148E-9 agidl = 0 bgidl = 2.3E9
+ cgidl = 0.5 egidl = 0.8 noia = 9E41
+ noib = 1E27 noic = 8E11 em = 4.1E7
+ af = 1 ef = 1.2 kf = 0
+ lintnoi = -3E-7 tnoia = 2.5E7 tnoib = 9.9E6
+ ntnoi = 1 rnoia = 0.912 rnoib = 0.26
+ xpart = 0 cgso = {2.392894381E-10/sw_func_tox_lv_ratio} cgdo = {2.392894381E-10/sw_func_tox_lv_ratio}
+ cgbo = {1E-14/sw_func_tox_lv_ratio} ckappas = 0.6 cf = 1E-14
+ clc = 1E-7 cle = 0.6 dlc = 1.21071E-8
+ dwc = 2.6E-8 vfbcv = -1 noff = 3.8661
+ voffcv = -0.16994 acde = 0.38008 moin = 23.81
+ cgsl = {2.310725E-11/sw_func_tox_lv_ratio} cgdl = {2.310725E-11/sw_func_tox_lv_ratio} ijthsrev = 0.1
+ ijthsfwd = 0.1 xjbvs = 1 bvs = 11.9
+ jss = 2.75E-3 jsws = 6E-10 cjs = {1.210E-03*sw_func_nsd_pw_cj}
+ mjs = 0.42197 mjsws = 1E-3 cjsws = {3.230311424E-11*sw_func_nsd_pw_cj}
+ cjswgs = {1.795291232E-10*sw_func_nsd_pw_cj} mjswgs = 0.8 pbs = 0.7477
+ pbsws = 0.1 pbswgs = 0.79644 xrcrg1 = 12
+ xrcrg2 = 1 rbpb = 50 rbpd = 50
+ rbps = 50 rbdb = 50 rbsb = 50
+ gbmin = 1E-12 tnom = 30 ute = -2.728772011666667
+ lute = 2.087495566594167E-7 wute = 2.216638084393335E-6 pute = -4.990059926062605E-13
+ kt1 = -0.9874280694 lkt1 = 1.0431523717593E-7 wkt1 = 2.678810021057867E-6
+ pkt1 = -4.103787081778183E-13 kt1l = 0 kt2 = -0.18195834168
+ lkt2 = 2.1358101945796E-8 wkt2 = 3.459564081993067E-7 pkt2 = -4.330130469812028E-14
+ ua1 = -5.818615500933333E-10 lua1 = 2.076285435242553E-16 wua1 = -5.59827440204854E-16
+ pua1 = -2.687278587551186E-22 ub1 = 3.831680610499996E-19 lub1 = -1.782357105377474E-25
+ wub1 = 3.391578918991267E-24 pub1 = -7.351384934137221E-32 uc1 = 7.131230292266665E-11
+ luc1 = -9.747080935509866E-18 wuc1 = 1.834316147919788E-16 puc1 = -3.540507207253452E-23
+ at = 2.935273537166666E5 lat = -0.029930442333614 wat = -0.863634922950067
+ pat = 1.203583353458449E-7 prt = 0 njs = 1.2928
+ xtis = 2 tpb = 1.2287E-3 tpbsw = 0
+ tpbswg = 0 tcj = 7.92E-4 tcjsw = 1E-5
+ tcjswg = 0 tvoff = 0 tvfbsdoff = 0
+ saref = 1.1E-6 sbref = 1.1E-6 wlod = 0
+ ku0 = -2.7E-8 kvsat = 0.2 kvth0 = 7.9E-9
+ tku0 = 0 llodku0 = 0 wlodku0 = 1
+ llodvth = 0 wlodvth = 1 lku0 = 0
+ wku0 = 0 pku0 = 0 lkvth0 = 0
+ wkvth0 = 3E-7 pkvth0 = 0 stk2 = 0
+ lodk2 = 1 steta0 = 0 lodeta0 = 1

.model nlowvt_model.25 nmos
+ level = 54 lmin = 8E-6 lmax = 2.02E-5 wmin = 1E-6
+ wmax = 3E-6 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 4.148E-9
+ toxm = 4.148E-9 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 9.999999999999999E22 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {2.6E-8+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {1.2025E-8-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = -1.33E-8 dwb = -1.08E-8 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = 0.431313765 wvth0 = -7.926479219999957E-9
+ vfb = 0 k1 = 0.49023394 wk1 = 4.078870487999991E-8
+ k2 = -0.045178254922 wk2 = -1.1596270717944E-8 k3 = 1.65
+ k3b = 1.6 w0 = 1E-7 lpe0 = 2.3802E-7
+ lpeb = -4.9152E-8 vbm = -3 dvtp0 = 0
+ dvtp1 = 0 dvt0 = 0.07665 dvt1 = 0.1252
+ dvt2 = -0.05637 dvt0w = 0 dvt1w = 5.3E6
+ dvt2w = -0.032 vfbsdoff = 0 u0 = 0.03333823146
+ wu0 = -2.020976224079999E-9 ua = -1.15871229168E-9 wua = 1.701070928726401E-16
+ ub = 2.55013008E-18 wub = -2.332459958400002E-25 uc = 9.11269848E-11
+ wuc = -6.520002511439999E-17 ud = 0 up = 0
+ lp = 1 eu = 1.67 vsat = 1.5520976E5
+ wvsat = 0.04298254752 a0 = 1.5719807236 wa0 = 3.306953680271999E-7
+ ags = 0.53432381 wags = 2.703876120000028E-9 b0 = 0
+ b1 = 0 keta = 0 a1 = 0
+ a2 = 0.38689047 rdsw = 103.65 rdswmin = 0
+ rdw = 0 rdwmin = 0 rsw = 0
+ rswmin = 0 prwb = 0 prwg = 0
+ wr = 1 voff = -0.11697059428 wvoff = 6.38620605744E-9
+ voffl = 0 minv = 0 nfactor = 1.16632463576
+ wnfactor = 4.9578993569952E-7 eta0 = 0.08 etab = -0.07
+ dsub = 0.56 cit = 2.63E-6 wcit = 6.98676E-12
+ cdsc = 3.8556E-37 cdscb = -1.1484E-4 cdscd = 4.7984E-6
+ pclm = 0.2 pdiblc1 = 0.39 pdiblc2 = 6.304997599999999E-3
+ wpdiblc2 = 1.1983690752E-9 pdiblcb = 0 drout = 3.4946
+ pscbe1 = 4.5E8 pscbe2 = 1E-8 pvag = 0
+ delta = 0.01 fprout = 0 pdits = 1.4427E-15
+ pditsl = 0 pditsd = 0 lambda = 0
+ vtl = 0 lc = 0 xn = 0
+ alpha0 = 3.7444087624E-5 walpha0 = 4.067725208447998E-12 alpha1 = 0
+ beta0 = 17.793363 aigbacc = 1 bigbacc = 0
+ cigbacc = 0 nigbacc = 1 aigbinv = 0.35
+ bigbinv = 0.03 cigbinv = 6E-3 eigbinv = 1.1
+ nigbinv = 3 aigc = 0.43 bigc = 0.054
+ cigc = 0.075 aigsd = 0.43 bigsd = 0.054
+ cigsd = 0.075 dlcig = 0 nigc = 1
+ poxedge = 1 pigcd = 1 ntox = 1
+ toxref = 4.148E-9 agidl = 0 bgidl = 2.3E9
+ cgidl = 0.5 egidl = 0.8 noia = 9E41
+ noib = 1E27 noic = 8E11 em = 4.1E7
+ af = 1 ef = 1.2 kf = 0
+ lintnoi = -3E-7 tnoia = 2.5E7 tnoib = 9.9E6
+ ntnoi = 1 rnoia = 0.912 rnoib = 0.26
+ xpart = 0 cgso = {2.392894381E-10/sw_func_tox_lv_ratio} cgdo = {2.392894381E-10/sw_func_tox_lv_ratio}
+ cgbo = {1E-14/sw_func_tox_lv_ratio} ckappas = 0.6 cf = 1E-14
+ clc = 1E-7 cle = 0.6 dlc = 1.21071E-8
+ dwc = 2.6E-8 vfbcv = -1 noff = 3.8661
+ voffcv = -0.16994 acde = 0.38008 moin = 23.81
+ cgsl = {2.310725E-11/sw_func_tox_lv_ratio} cgdl = {2.310725E-11/sw_func_tox_lv_ratio} ijthsrev = 0.1
+ ijthsfwd = 0.1 xjbvs = 1 bvs = 11.9
+ jss = 2.75E-3 jsws = 6E-10 cjs = {1.210E-03*sw_func_nsd_pw_cj}
+ mjs = 0.42197 mjsws = 1E-3 cjsws = {3.230311424E-11*sw_func_nsd_pw_cj}
+ cjswgs = {1.795291232E-10*sw_func_nsd_pw_cj} mjswgs = 0.8 pbs = 0.7477
+ pbsws = 0.1 pbswgs = 0.79644 xrcrg1 = 12
+ xrcrg2 = 1 rbpb = 50 rbpd = 50
+ rbps = 50 rbdb = 50 rbsb = 50
+ gbmin = 1E-12 tnom = 30 ute = -1.2990148
+ wute = 1.120676303999998E-7 kt1 = -0.25493258 wkt1 = -2.557154159999997E-9
+ kt1l = 0 kt2 = -0.034029184 wkt2 = -2.213405568000003E-9
+ ua1 = 2.1423962E-9 wua1 = -1.694987976E-16 ub1 = -2.3838598E-18
+ wub1 = 8.701310904E-25 uc1 = -9.907576E-11 wuc1 = 1.5404408448E-16
+ at = 4.418385E5 wat = -0.363660858 prt = 0
+ njs = 1.2928 xtis = 2 tpb = 1.2287E-3
+ tpbsw = 0 tpbswg = 0 tcj = 7.92E-4
+ tcjsw = 1E-5 tcjswg = 0 tvoff = 0
+ tvfbsdoff = 0 saref = 3E-6 sbref = 3E-6
+ wlod = 0 ku0 = -2.7E-8 kvsat = 0.2
+ kvth0 = 7.9E-9 tku0 = 0 llodku0 = 0
+ wlodku0 = 1 llodvth = 0 wlodvth = 1
+ lku0 = 0 wku0 = 0 pku0 = 0
+ lkvth0 = 0 wkvth0 = 3E-7 pkvth0 = 0
+ stk2 = 0 lodk2 = 1 steta0 = 0
+ lodeta0 = 1

.model nlowvt_model.26 nmos
+ level = 54 lmin = 4E-6 lmax = 8E-6 wmin = 1E-6
+ wmax = 3E-6 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 4.148E-9
+ toxm = 4.148E-9 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 9.999999999999999E22 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {2.6E-8+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {1.2025E-8-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = -1.33E-8 dwb = -1.08E-8 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = 0.431313765 wvth0 = -7.926479219999957E-9
+ vfb = 0 k1 = 0.49023394 wk1 = 4.078870487999991E-8
+ k2 = -0.045178254922 wk2 = -1.1596270717944E-8 k3 = 1.65
+ k3b = 1.6 w0 = 1E-7 lpe0 = 2.3802E-7
+ lpeb = -4.9152E-8 vbm = -3 dvtp0 = 0
+ dvtp1 = 0 dvt0 = 0.07665 dvt1 = 0.1252
+ dvt2 = -0.05637 dvt0w = 0 dvt1w = 5.3E6
+ dvt2w = -0.032 vfbsdoff = 0 u0 = 0.03333823146
+ wu0 = -2.020976224079999E-9 ua = -1.15871229168E-9 wua = 1.701070928726401E-16
+ ub = 2.55013008E-18 wub = -2.332459958400002E-25 uc = 9.11269848E-11
+ wuc = -6.520002511439999E-17 ud = 0 up = 0
+ lp = 1 eu = 1.67 vsat = 1.5520976E5
+ wvsat = 0.04298254752 a0 = 1.5719807236 wa0 = 3.306953680271999E-7
+ ags = 0.53432381 wags = 2.703876120000028E-9 b0 = 0
+ b1 = 0 keta = 0 a1 = 0
+ a2 = 0.38689047 rdsw = 103.65 rdswmin = 0
+ rdw = 0 rdwmin = 0 rsw = 0
+ rswmin = 0 prwb = 0 prwg = 0
+ wr = 1 voff = -0.11697059428 wvoff = 6.38620605744E-9
+ voffl = 0 minv = 0 nfactor = 1.16632463576
+ wnfactor = 4.9578993569952E-7 eta0 = 0.08 etab = -0.07
+ dsub = 0.56 cit = 2.63E-6 wcit = 6.98676E-12
+ cdsc = 3.8556E-37 cdscb = -1.1484E-4 cdscd = 4.7984E-6
+ pclm = 0.2 pdiblc1 = 0.39 pdiblc2 = 6.304997599999999E-3
+ wpdiblc2 = 1.1983690752E-9 pdiblcb = 0 drout = 3.4946
+ pscbe1 = 4.5E8 pscbe2 = 1E-8 pvag = 0
+ delta = 0.01 fprout = 0 pdits = 1.4427E-15
+ pditsl = 0 pditsd = 0 lambda = 0
+ vtl = 0 lc = 0 xn = 0
+ alpha0 = 3.7444087624E-5 walpha0 = 4.067725208447998E-12 alpha1 = 0
+ beta0 = 17.793363 aigbacc = 1 bigbacc = 0
+ cigbacc = 0 nigbacc = 1 aigbinv = 0.35
+ bigbinv = 0.03 cigbinv = 6E-3 eigbinv = 1.1
+ nigbinv = 3 aigc = 0.43 bigc = 0.054
+ cigc = 0.075 aigsd = 0.43 bigsd = 0.054
+ cigsd = 0.075 dlcig = 0 nigc = 1
+ poxedge = 1 pigcd = 1 ntox = 1
+ toxref = 4.148E-9 agidl = 0 bgidl = 2.3E9
+ cgidl = 0.5 egidl = 0.8 noia = 9E41
+ noib = 1E27 noic = 8E11 em = 4.1E7
+ af = 1 ef = 1.2 kf = 0
+ lintnoi = -3E-7 tnoia = 2.5E7 tnoib = 9.9E6
+ ntnoi = 1 rnoia = 0.912 rnoib = 0.26
+ xpart = 0 cgso = {2.392894381E-10/sw_func_tox_lv_ratio} cgdo = {2.392894381E-10/sw_func_tox_lv_ratio}
+ cgbo = {1E-14/sw_func_tox_lv_ratio} ckappas = 0.6 cf = 1E-14
+ clc = 1E-7 cle = 0.6 dlc = 1.21071E-8
+ dwc = 2.6E-8 vfbcv = -1 noff = 3.8661
+ voffcv = -0.16994 acde = 0.38008 moin = 23.81
+ cgsl = {2.310725E-11/sw_func_tox_lv_ratio} cgdl = {2.310725E-11/sw_func_tox_lv_ratio} ijthsrev = 0.1
+ ijthsfwd = 0.1 xjbvs = 1 bvs = 11.9
+ jss = 2.75E-3 jsws = 6E-10 cjs = {1.210E-03*sw_func_nsd_pw_cj}
+ mjs = 0.42197 mjsws = 1E-3 cjsws = {3.230311424E-11*sw_func_nsd_pw_cj}
+ cjswgs = {1.795291232E-10*sw_func_nsd_pw_cj} mjswgs = 0.8 pbs = 0.7477
+ pbsws = 0.1 pbswgs = 0.79644 xrcrg1 = 12
+ xrcrg2 = 1 rbpb = 50 rbpd = 50
+ rbps = 50 rbdb = 50 rbsb = 50
+ gbmin = 1E-12 tnom = 30 ute = -1.2990148
+ wute = 1.120676303999998E-7 kt1 = -0.25493258 wkt1 = -2.557154159999997E-9
+ kt1l = 0 kt2 = -0.034029184 wkt2 = -2.213405568000003E-9
+ ua1 = 2.1423962E-9 wua1 = -1.694987976E-16 ub1 = -2.3838598E-18
+ wub1 = 8.701310904E-25 uc1 = -9.907576E-11 wuc1 = 1.5404408448E-16
+ at = 4.418385E5 wat = -0.363660858 prt = 0
+ njs = 1.2928 xtis = 2 tpb = 1.2287E-3
+ tpbsw = 0 tpbswg = 0 tcj = 7.92E-4
+ tcjsw = 1E-5 tcjswg = 0 tvoff = 0
+ tvfbsdoff = 0 saref = 3E-6 sbref = 3E-6
+ wlod = 0 ku0 = -2.7E-8 kvsat = 0.2
+ kvth0 = 7.9E-9 tku0 = 0 llodku0 = 0
+ wlodku0 = 1 llodvth = 0 wlodvth = 1
+ lku0 = 0 wku0 = 0 pku0 = 0
+ lkvth0 = 0 wkvth0 = 3E-7 pkvth0 = 0
+ stk2 = 0 lodk2 = 1 steta0 = 0
+ lodeta0 = 1

.model nlowvt_model.27 nmos
+ level = 54 lmin = 2E-6 lmax = 4E-6 wmin = 1E-6
+ wmax = 3E-6 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 4.148E-9
+ toxm = 4.148E-9 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 9.999999999999999E22 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {2.6E-8+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {1.2025E-8-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = -1.33E-8 dwb = -1.08E-8 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = 0.426562078094835 lvth0 = 1.889246955059097E-8
+ wvth0 = -1.372326575351347E-8 pvth0 = 2.304773341792305E-14 vfb = 0
+ k1 = 0.544648876189 lk1 = -2.163510655406545E-7 wk1 = 5.975744597182788E-8
+ pk1 = -7.541876614405341E-14 k2 = -0.072613436357313 lk2 = 1.090809096277326E-7
+ wk2 = -1.328571322193972E-8 pk2 = 6.717138923761784E-15 k3 = 1.65
+ k3b = 1.6 w0 = 1E-7 lpe0 = 2.3802E-7
+ lpeb = -4.9152E-8 vbm = -3 dvtp0 = 0
+ dvtp1 = 0 dvt0 = 0.07665 dvt1 = 0.1252
+ dvt2 = -0.05637 dvt0w = 0 dvt1w = 5.3E6
+ dvt2w = -0.032 vfbsdoff = 0 u0 = 0.034060244617494
+ lu0 = -2.870688213538278E-9 wu0 = -2.918277749556314E-9 pu0 = 3.567626000217552E-15
+ ua = -1.023713958020897E-9 lua = -5.367466247119121E-16 wua = 1.637694211082412E-16
+ pua = 2.519826605166185E-23 ub = 2.4366531091335E-18 lub = 4.51178762316661E-25
+ wub = -2.896966379975584E-25 pub = 2.244449306863437E-31 uc = 7.577744241557997E-11
+ luc = 6.102901304333477E-17 wuc = -7.791722688409372E-17 puc = 5.056295837621378E-23
+ ud = 0 up = 0 lp = 1
+ eu = 1.67 vsat = 2.7304558764875E5 lvsat = -0.468509358940048
+ wvsat = 0.079118413464585 pvsat = -1.436743962023728E-7 a0 = 1.30855970935696
+ la0 = 1.047348781579615E-6 wa0 = 6.449132544877518E-7 pa0 = -1.249314605672831E-12
+ ags = -0.8435163683248 lags = 5.47822365701049E-6 wags = 4.525308664717105E-7
+ pags = -1.788489622288883E-12 b0 = 0 b1 = 0
+ keta = 0.281834609337 lketa = -1.120560314993445E-6 wketa = -9.743913728247601E-8
+ pketa = 3.874131378782604E-13 a1 = 0 a2 = 0.38689047
+ rdsw = 103.65 rdswmin = 0 rdw = 0
+ rdwmin = 0 rsw = 0 rswmin = 0
+ prwb = 0 prwg = 0 wr = 1
+ voff = -0.11564535387882 lvoff = -5.269089573073569E-9 wvoff = 1.150408008682489E-8
+ pvoff = -2.034841124713286E-14 voffl = 0 minv = 0
+ nfactor = 1.025218886794988 lnfactor = 5.610294025974395E-7 wnfactor = 9.705815012086405E-7
+ pnfactor = -1.887747524885987E-12 eta0 = 0.1585440125 leta0 = -3.122870664993751E-7
+ etab = -0.138675665134425 letab = 2.730510107912152E-7 wetab = 1.080969743442647E-11
+ petab = -4.297881651440792E-17 dsub = 0.800343584265283 ldsub = -9.555940738595502E-7
+ wdsub = -8.00905392844118E-8 pdsub = 3.18435979667857E-13 cit = 2.63E-6
+ wcit = 6.98676E-12 cdsc = 3.8556E-37 cdscb = -1.1484E-4
+ cdscd = 4.7984E-6 pclm = 0.2398203126155 lpclm = -1.583235719435972E-7
+ wpclm = -7.0090464718494E-8 ppclm = 2.786761831974962E-13 pdiblc1 = 0.39
+ pdiblc2 = 6.410177616095001E-3 lpdiblc2 = -4.181904849929193E-10 wpdiblc2 = -2.815300573728063E-9
+ ppdiblc2 = 1.595814984065553E-14 pdiblcb = 0 drout = 3.4946
+ pscbe1 = 4.5E8 pscbe2 = 1E-8 pvag = 0
+ delta = 0.01 fprout = 0 pdits = 1.4427E-15
+ pditsl = 0 pditsd = 0 lambda = 0
+ vtl = 0 lc = 0 xn = 0
+ alpha0 = -7.409723927919266E-5 lalpha0 = 4.434827387007488E-10 walpha0 = 3.235211168889172E-11
+ palpha0 = -1.124573064269202E-16 alpha1 = 0 beta0 = 14.038366508569252
+ lbeta0 = 1.494366743367018E-5 wbeta0 = 3.772887393147458E-7 pbeta0 = -1.51334286169914E-12
+ aigbacc = 1 bigbacc = 0 cigbacc = 0
+ nigbacc = 1 aigbinv = 0.35 bigbinv = 0.03
+ cigbinv = 6E-3 eigbinv = 1.1 nigbinv = 3
+ aigc = 0.43 bigc = 0.054 cigc = 0.075
+ aigsd = 0.43 bigsd = 0.054 cigsd = 0.075
+ dlcig = 0 nigc = 1 poxedge = 1
+ pigcd = 1 ntox = 1 toxref = 4.148E-9
+ agidl = 0 bgidl = 2.3E9 cgidl = 0.5
+ egidl = 0.8 noia = 9E41 noib = 1E27
+ noic = 8E11 em = 4.1E7 af = 1
+ ef = 1.2 kf = 0 lintnoi = -3E-7
+ tnoia = 2.5E7 tnoib = 9.9E6 ntnoi = 1
+ rnoia = 0.912 rnoib = 0.26 xpart = 0
+ cgso = {2.392894381E-10/sw_func_tox_lv_ratio} cgdo = {2.392894381E-10/sw_func_tox_lv_ratio} cgbo = {1E-14/sw_func_tox_lv_ratio}
+ ckappas = 0.6 cf = 1E-14 clc = 1E-7
+ cle = 0.6 dlc = 1.21071E-8 dwc = 2.6E-8
+ vfbcv = -1 noff = 3.8661 voffcv = -0.16994
+ acde = 0.38008 moin = 23.81 cgsl = {2.310725E-11/sw_func_tox_lv_ratio}
+ cgdl = {2.310725E-11/sw_func_tox_lv_ratio} ijthsrev = 0.1 ijthsfwd = 0.1
+ xjbvs = 1 bvs = 11.9 jss = 2.75E-3
+ jsws = 6E-10 cjs = {1.210E-03*sw_func_nsd_pw_cj} mjs = 0.42197
+ mjsws = 1E-3 cjsws = {3.230311424E-11*sw_func_nsd_pw_cj} cjswgs = {1.795291232E-10*sw_func_nsd_pw_cj}
+ mjswgs = 0.8 pbs = 0.7477 pbsws = 0.1
+ pbswgs = 0.79644 xrcrg1 = 12 xrcrg2 = 1
+ rbpb = 50 rbpd = 50 rbps = 50
+ rbdb = 50 rbsb = 50 gbmin = 1E-12
+ tnom = 30 ute = -1.34423481094 lute = 1.797925024968926E-7
+ wute = 9.770992244111949E-8 pute = 5.708552895910998E-14 kt1 = -0.2634400524845
+ lkt1 = 3.382528522474776E-8 wkt1 = 1.570750702230596E-8 pkt1 = -7.261937962778937E-14
+ kt1l = 0 kt2 = -0.03223380223885 lkt2 = -7.138348113244364E-9
+ wkt2 = -3.236392260070211E-9 pkt2 = 4.067343938336544E-15 ua1 = 1.97185788335E-9
+ lua1 = 6.780518200845672E-16 wua1 = -8.528531822579979E-17 pua1 = -3.348285833178512E-22
+ ub1 = -1.985903667595E-18 lub1 = -1.58225368463566E-24 wub1 = 8.9401458537006E-25
+ pub1 = -9.49595818262106E-32 uc1 = -1.23373526521615E-10 luc1 = 9.66067048016152E-17
+ wuc1 = 2.450831353849211E-16 puc1 = -3.619667144454208E-22 at = 8.391688786792503E5
+ lat = -1.579765719109764 wat = -0.731846331470529 pat = 1.46388703324515E-6
+ prt = 0 njs = 1.2928 xtis = 2
+ tpb = 1.2287E-3 tpbsw = 0 tpbswg = 0
+ tcj = 7.92E-4 tcjsw = 1E-5 tcjswg = 0
+ tvoff = 0 tvfbsdoff = 0 saref = 3E-6
+ sbref = 3E-6 wlod = 0 ku0 = -2.7E-8
+ kvsat = 0.2 kvth0 = 7.9E-9 tku0 = 0
+ llodku0 = 0 wlodku0 = 1 llodvth = 0
+ wlodvth = 1 lku0 = 0 wku0 = 0
+ pku0 = 0 lkvth0 = 0 wkvth0 = 3E-7
+ pkvth0 = 0 stk2 = 0 lodk2 = 1
+ steta0 = 0 lodeta0 = 1

.model nlowvt_model.28 nmos
+ level = 54 lmin = 1E-6 lmax = 2E-6 wmin = 1E-6
+ wmax = 3E-6 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 4.148E-9
+ toxm = 4.148E-9 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 9.999999999999999E22 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {2.6E-8+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {1.2025E-8-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = -1.33E-8 dwb = -1.08E-8 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = 0.435697877817309 lvth0 = 8.405860889682165E-10
+ wvth0 = -5.994948864749011E-9 pvth0 = 7.776965661568916E-15 vfb = 0
+ k1 = 0.441796029293 lk1 = -1.31189827165033E-8 wk1 = 1.571134450023605E-8
+ pk1 = 1.161412805873862E-14 k2 = -0.01392863337349 lk2 = -6.877326828152431E-9
+ wk2 = -8.824862133831479E-9 pk2 = -2.097279783785694E-15 k3 = 1.65
+ k3b = 1.6 w0 = 1E-7 lpe0 = 2.3802E-7
+ lpeb = -4.9152E-8 vbm = -3 dvtp0 = 0
+ dvtp1 = 0 dvt0 = 0.07665 dvt1 = 0.1252
+ dvt2 = -0.05637 dvt0w = 0 dvt1w = 5.3E6
+ dvt2w = -0.032 vfbsdoff = 0 u0 = 0.035918173255615
+ lu0 = -6.541862306034241E-9 wu0 = 2.200107917818074E-10 pu0 = -2.633475243039509E-15
+ ua = -1.116781612163862E-9 lua = -3.528495935081202E-16 wua = 3.780624313715588E-16
+ pua = -3.982340075781406E-22 ub = 2.667103533068E-18 lub = -4.179752856714329E-27
+ wub = -2.968815903704638E-25 pub = 2.386420373275861E-31 uc = 1.255958958374E-10
+ luc = -3.740975999551056E-17 wuc = -6.386259869465522E-17 puc = 2.279171580529277E-23
+ ud = 0 up = 0 lp = 1
+ eu = 1.67 vsat = -2.500485490799998E3 lvsat = 0.075955904280046
+ wvsat = 4.546709806478401E-3 pvsat = 3.675561640863004E-9 a0 = 2.0849995442401
+ la0 = -4.868575101577254E-7 wa0 = 1.238432992461853E-7 pa0 = -2.197064276132578E-13
+ ags = 1.6265133855182 lags = 5.975683649044128E-7 wags = -4.108593203272532E-7
+ pags = -8.247378268347039E-14 b0 = 0 b1 = 0
+ keta = -0.348937225292 lketa = 1.258132916417273E-7 wketa = 9.540666434481593E-8
+ pketa = 6.359476152812901E-15 a1 = 0 a2 = 0.38689047
+ rdsw = 103.65 rdswmin = 0 rdw = 0
+ rdwmin = 0 rsw = 0 rswmin = 0
+ prwb = 0 prwg = 0 wr = 1
+ voff = -0.120031162167445 lvoff = 3.397048314835952E-9 wvoff = 1.087599224989856E-9
+ pvoff = 2.340341118100805E-16 voffl = 0 minv = 0
+ nfactor = 0.814253125507248 lnfactor = 9.778871986139493E-7 wnfactor = -7.643669107078897E-8
+ pnfactor = 1.811080721485515E-13 eta0 = 5.18411862801E-4 leta0 = -3.638092030163599E-11
+ weta0 = 4.408989797665201E-11 peta0 = -8.711943390696552E-17 etab = -5.03400784399E-4
+ letab = 2.952504878220398E-11 wetab = -2.276494124374802E-11 petab = 2.336299078173188E-17
+ dsub = -0.238858339241776 ldsub = 1.097816966894222E-6 wdsub = 4.500279996800494E-7
+ pdsub = -7.290517473989701E-13 cit = 3.169984999999997E-7 lcit = 4.570375313924999E-12
+ wcit = 1.3805488422E-11 pcit = -1.34734664254509E-17 cdsc = 3.8556E-37
+ cdscb = -1.1484E-4 cdscd = 4.7984E-6 pclm = 0.284056561333
+ lpclm = -2.457321875969414E-7 wpclm = -2.603239457768406E-8 ppclm = 1.916196395027628E-13
+ pdiblc1 = 0.39 pdiblc2 = 1.584281503000081E-5 lpdiblc2 = 1.221669536517147E-8
+ wpdiblc2 = 8.39736924435156E-9 ppdiblc2 = -6.197525086378905E-15 pdiblcb = 0
+ drout = 3.4946 pscbe1 = 4.5E8 pscbe2 = 1E-8
+ pvag = 0 delta = 0.01 fprout = 0
+ pdits = 1.4427E-15 pditsl = 0 pditsd = 0
+ lambda = 0 vtl = 0 lc = 0
+ xn = 0 alpha0 = 2.508406437580834E-4 lalpha0 = -1.985782712867569E-10
+ walpha0 = -4.824410741611072E-11 palpha0 = 4.679679271360937E-17 alpha1 = 0
+ beta0 = 22.352715437401 lbeta0 = -1.485070332254902E-6 wbeta0 = -7.140775948797478E-7
+ pbeta0 = 6.431424463524706E-13 aigbacc = 1 bigbacc = 0
+ cigbacc = 0 nigbacc = 1 aigbinv = 0.35
+ bigbinv = 0.03 cigbinv = 6E-3 eigbinv = 1.1
+ nigbinv = 3 aigc = 0.43 bigc = 0.054
+ cigc = 0.075 aigsd = 0.43 bigsd = 0.054
+ cigsd = 0.075 dlcig = 0 nigc = 1
+ poxedge = 1 pigcd = 1 ntox = 1
+ toxref = 4.148E-9 agidl = 0 bgidl = 2.3E9
+ cgidl = 0.5 egidl = 0.8 noia = 9E41
+ noib = 1E27 noic = 8E11 em = 4.1E7
+ af = 1 ef = 1.2 kf = 0
+ lintnoi = -3E-7 tnoia = 2.5E7 tnoib = 9.9E6
+ ntnoi = 1 rnoia = 0.912 rnoib = 0.26
+ xpart = 0 cgso = {2.392894381E-10/sw_func_tox_lv_ratio} cgdo = {2.392894381E-10/sw_func_tox_lv_ratio}
+ cgbo = {1E-14/sw_func_tox_lv_ratio} ckappas = 0.6 cf = 1E-14
+ clc = 1E-7 cle = 0.6 dlc = 1.21071E-8
+ dwc = 2.6E-8 vfbcv = -1 noff = 3.8661
+ voffcv = -0.16994 acde = 0.38008 moin = 23.81
+ cgsl = {2.310725E-11/sw_func_tox_lv_ratio} cgdl = {2.310725E-11/sw_func_tox_lv_ratio} ijthsrev = 0.1
+ ijthsfwd = 0.1 xjbvs = 1 bvs = 11.9
+ jss = 2.75E-3 jsws = 6E-10 cjs = {1.210E-03*sw_func_nsd_pw_cj}
+ mjs = 0.42197 mjsws = 1E-3 cjsws = {3.230311424E-11*sw_func_nsd_pw_cj}
+ cjswgs = {1.795291232E-10*sw_func_nsd_pw_cj} mjswgs = 0.8 pbs = 0.7477
+ pbsws = 0.1 pbswgs = 0.79644 xrcrg1 = 12
+ xrcrg2 = 1 rbpb = 50 rbpd = 50
+ rbps = 50 rbdb = 50 rbsb = 50
+ gbmin = 1E-12 tnom = 30 ute = -1.39045594316
+ lute = 2.711231487070017E-7 wute = 2.318812580356799E-7 pute = -2.080303216089617E-13
+ kt1 = -0.229914591284 lkt1 = -3.241934983438008E-8 wkt1 = -3.566347485676788E-8
+ pkt1 = 2.888711201616659E-14 kt1l = 0 kt2 = -0.0512034811769
+ lkt2 = 3.034478898439556E-8 wkt2 = 8.076953070121421E-11 pkt2 = -2.487201902138255E-15
+ ua1 = 1.61399917349E-9 lua1 = 1.385162737832435E-15 wua1 = 4.567288539514796E-16
+ pua1 = -1.405821486831546E-21 ub1 = -1.90303076139E-18 lub1 = -1.746006403651429E-24
+ wub1 = -1.4780457942228E-25 pub1 = 1.963622996845214E-30 uc1 = -4.394409656867002E-11
+ luc1 = -6.03418773139065E-17 wuc1 = 7.066434908723916E-17 puc1 = -1.732391366051626E-23
+ at = 3.768967792500002E3 lat = 0.07094273480691 wat = 0.01585875570411
+ pat = -1.354083375757815E-8 prt = 0 njs = 1.2928
+ xtis = 2 tpb = 1.2287E-3 tpbsw = 0
+ tpbswg = 0 tcj = 7.92E-4 tcjsw = 1E-5
+ tcjswg = 0 tvoff = 0 tvfbsdoff = 0
+ saref = 3E-6 sbref = 3E-6 wlod = 0
+ ku0 = -2.7E-8 kvsat = 0.2 kvth0 = 7.9E-9
+ tku0 = 0 llodku0 = 0 wlodku0 = 1
+ llodvth = 0 wlodvth = 1 lku0 = 0
+ wku0 = 0 pku0 = 0 lkvth0 = 0
+ wkvth0 = 3E-7 pkvth0 = 0 stk2 = 0
+ lodk2 = 1 steta0 = 0 lodeta0 = 1

.model nlowvt_model.29 nmos
+ level = 54 lmin = 5E-7 lmax = 1E-6 wmin = 1E-6
+ wmax = 3E-6 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 4.148E-9
+ toxm = 4.148E-9 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 9.999999999999999E22 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {2.6E-8+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {1.2025E-8-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = -1.33E-8 dwb = -1.08E-8 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = 0.444062643187062 lvth0 = -7.323006673642111E-9
+ wvth0 = 2.68293210098532E-9 pvth0 = -6.922122669395036E-16 vfb = 0
+ k1 = 0.444861876332 lk1 = -1.611109613421537E-8 wk1 = -1.944021254735951E-9
+ pk1 = 2.884488226730355E-14 k2 = -0.021767612643805 lk2 = 7.731249907114908E-10
+ wk2 = -1.290177082346467E-9 pk2 = -9.45075565978249E-15 k3 = 1.65
+ k3b = 1.6 w0 = 1E-7 lpe0 = 2.3802E-7
+ lpeb = -4.9152E-8 vbm = -3 dvtp0 = 0
+ dvtp1 = 0 dvt0 = 0.07665 dvt1 = 0.1252
+ dvt2 = -0.05637 dvt0w = 0 dvt1w = 5.3E6
+ dvt2w = -0.032 vfbsdoff = 0 u0 = 0.027351692126439
+ lu0 = 1.818594951985262E-9 wu0 = 2.926352457361234E-9 pu0 = -5.27472939156175E-15
+ ua = -1.954136517320322E-9 lua = 4.643669261793273E-16 wua = 7.247943112586693E-16
+ pua = -7.36626985753966E-22 ub = 3.311994286502E-18 lub = -6.335608836706269E-25
+ wub = -7.09673751319896E-25 pub = 6.415065468061845E-31 uc = 1.280887001497826E-10
+ luc = -3.984261236418032E-17 wuc = -9.024443704475909E-17 puc = 4.853907094307664E-23
+ ud = 0 up = 0 lp = 1
+ eu = 1.67 vsat = -1.276653505661998E4 lvsat = 0.085975055353808
+ wvsat = 0.012872165762436 pvsat = -4.449667099353557E-9 a0 = 1.0027629971188
+ la0 = 5.693512480053072E-7 wa0 = 9.040447169617774E-7 pa0 = -9.811440012327898E-13
+ ags = 3.3381908499998 lags = -1.072943256556405E-6 wags = -1.932017060638106E-7
+ pags = -2.948967313238772E-13 b0 = 0 b1 = 0
+ keta = -0.412482366837846 lketa = 1.878301725333954E-7 wketa = 1.828446447502776E-7
+ pketa = -7.897562082389746E-14 a1 = 0 a2 = 0.38689047
+ rdsw = 103.65 rdswmin = 0 rdw = 0
+ rdwmin = 0 rsw = 0 rswmin = 0
+ prwb = 0 prwg = 0 wr = 1
+ voff = -0.12697698918715 lvoff = 1.017582819471705E-8 wvoff = 1.81406947153542E-8
+ pvoff = -1.6408934432011E-14 voffl = 0 minv = 0
+ nfactor = 1.104843260815356 lnfactor = 6.942857560600014E-7 wnfactor = 4.318497725189629E-7
+ pnfactor = -3.149541019918668E-13 eta0 = 2.147920770653582E-3 leta0 = -1.626700138920362E-9
+ weta0 = -3.679767982914753E-9 peta0 = 3.547179664949001E-15 etab = -8.404806148316381E-4
+ letab = 3.584981092929371E-10 wetab = 3.635294256839287E-11 petab = -3.433310792472702E-17
+ dsub = 0.777506341422422 ldsub = 1.058958567999982E-7 wdsub = -5.796938422224519E-7
+ pdsub = 2.759052842057759E-13 cit = 5E-6 cdsc = 3.8556E-37
+ cdscb = -1.1484E-4 cdscd = 4.7984E-6 pclm = -0.203163899708
+ lpclm = 2.297706213560226E-7 wpclm = 2.91591369407184E-7 ppclm = -1.183652729582692E-13
+ pdiblc1 = 0.39 pdiblc2 = 0.01246240729876 lpdiblc2 = 6.947075727518027E-11
+ wpdiblc2 = 8.74490445765552E-9 ppdiblc2 = -6.536702077802904E-15 pdiblcb = 0
+ drout = 3.4946 pscbe1 = 4.5E8 pscbe2 = 1E-8
+ pvag = 0 delta = 0.01 fprout = 0
+ pdits = 1.4427E-15 pditsl = 0 pditsd = 0
+ lambda = 0 vtl = 0 lc = 0
+ xn = 0 alpha0 = 2.162008659521218E-6 lalpha0 = 4.411964263768487E-11
+ walpha0 = -4.206475273024288E-11 palpha0 = 4.076605150793666E-17 alpha1 = 0
+ beta0 = 18.299816647158405 lbeta0 = 2.470356242082357E-6 wbeta0 = -8.242581225037668E-7
+ pbeta0 = 7.506731322871318E-13 aigbacc = 1 bigbacc = 0
+ cigbacc = 0 nigbacc = 1 aigbinv = 0.35
+ bigbinv = 0.03 cigbinv = 6E-3 eigbinv = 1.1
+ nigbinv = 3 aigc = 0.43 bigc = 0.054
+ cigc = 0.075 aigsd = 0.43 bigsd = 0.054
+ cigsd = 0.075 dlcig = 0 nigc = 1
+ poxedge = 1 pigcd = 1 ntox = 1
+ toxref = 4.148E-9 agidl = 0 bgidl = 2.3E9
+ cgidl = 0.5 egidl = 0.8 noia = 9E41
+ noib = 1E27 noic = 8E11 em = 4.1E7
+ af = 1 ef = 1.2 kf = 0
+ lintnoi = -3E-7 tnoia = 2.5E7 tnoib = 9.9E6
+ ntnoi = 1 rnoia = 0.912 rnoib = 0.26
+ xpart = 0 cgso = {2.392894381E-10/sw_func_tox_lv_ratio} cgdo = {2.392894381E-10/sw_func_tox_lv_ratio}
+ cgbo = {1E-14/sw_func_tox_lv_ratio} ckappas = 0.6 cf = 1E-14
+ clc = 1E-7 cle = 0.6 dlc = 1.21071E-8
+ dwc = 2.6E-8 vfbcv = -1 noff = 3.8661
+ voffcv = -0.16994 acde = 0.38008 moin = 23.81
+ cgsl = {2.310725E-11/sw_func_tox_lv_ratio} cgdl = {2.310725E-11/sw_func_tox_lv_ratio} ijthsrev = 0.1
+ ijthsfwd = 0.1 xjbvs = 1 bvs = 11.9
+ jss = 2.75E-3 jsws = 6E-10 cjs = {1.210E-03*sw_func_nsd_pw_cj}
+ mjs = 0.42197 mjsws = 1E-3 cjsws = {3.230311424E-11*sw_func_nsd_pw_cj}
+ cjswgs = {1.795291232E-10*sw_func_nsd_pw_cj} mjswgs = 0.8 pbs = 0.7477
+ pbsws = 0.1 pbswgs = 0.79644 xrcrg1 = 12
+ xrcrg2 = 1 rbpb = 50 rbpd = 50
+ rbps = 50 rbdb = 50 rbsb = 50
+ gbmin = 1E-12 tnom = 30 ute = -0.51727832018
+ lute = -5.810545524403289E-7 wute = -5.129321889093598E-7 pute = 5.188703619370498E-13
+ kt1 = -0.273206835776 lkt1 = 9.83171617758717E-9 wkt1 = 4.523401695647941E-9
+ pkt1 = -1.033327015516362E-14 kt1l = 0 kt2 = -0.0204380516654
+ lkt2 = 3.192680526471342E-10 wkt2 = 9.648515878399203E-9 pkt2 = -1.18248439501741E-14
+ ua1 = 6.165976834958001E-9 lua1 = -3.05733986087726E-15 wua1 = -3.471003317900184E-15
+ pua1 = 2.427448726287085E-21 ub1 = -7.69693020612E-18 lub1 = 3.908549759432813E-24
+ wub1 = 5.269630115201759E-24 pub1 = -3.323522393373116E-30 uc1 = -2.117399909437999E-10
+ luc1 = 1.034185258015016E-16 wuc1 = 1.188525271135224E-16 puc1 = -6.435316600526736E-23
+ at = 8.513982966900001E4 lat = -8.47115784146055E-3 wat = -8.809841137812E-3
+ pat = 1.053448333029562E-8 prt = 0 njs = 1.2928
+ xtis = 2 tpb = 1.2287E-3 tpbsw = 0
+ tpbswg = 0 tcj = 7.92E-4 tcjsw = 1E-5
+ tcjswg = 0 tvoff = 0 tvfbsdoff = 0
+ saref = 2.74E-6 sbref = 2.74E-6 wlod = 0
+ ku0 = -2.7E-8 kvsat = 0.2 kvth0 = 7.9E-9
+ tku0 = 0 llodku0 = 0 wlodku0 = 1
+ llodvth = 0 wlodvth = 1 lku0 = 0
+ wku0 = 0 pku0 = 0 lkvth0 = 0
+ wkvth0 = 3E-7 pkvth0 = 0 stk2 = 0
+ lodk2 = 1 steta0 = 0 lodeta0 = 1

.model nlowvt_model.30 nmos
+ level = 54 lmin = 2.5E-7 lmax = 5E-7 wmin = 1E-6
+ wmax = 3E-6 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 4.148E-9
+ toxm = 4.148E-9 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 9.999999999999999E22 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {2.6E-8+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {1.2025E-8-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = -1.33E-8 dwb = -1.08E-8 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = 0.495732629876516 lvth0 = -3.191533683848779E-8
+ wvth0 = -1.29637423017267E-10 pvth0 = 6.464301980095274E-16 vfb = 0
+ k1 = 0.253459673991752 lk1 = 7.498678206962564E-8 wk1 = 9.867482676781907E-8
+ pk1 = -1.904465844903151E-14 k2 = 0.030027345789938 lk2 = -2.387868547582849E-8
+ wk2 = -3.965639106104044E-8 pk2 = 8.809643883376904E-15 k3 = 1.65
+ k3b = 1.6 w0 = 1E-7 lpe0 = 2.3802E-7
+ lpeb = -4.9152E-8 vbm = -3 dvtp0 = 0
+ dvtp1 = 0 dvt0 = 0.07665 dvt1 = 0.1252
+ dvt2 = -0.05637 dvt0w = 0 dvt1w = 5.3E6
+ dvt2w = -0.032 vfbsdoff = 0 u0 = 0.040037742454812
+ lu0 = -4.219330701803961E-9 wu0 = -1.255264745337815E-8 pu0 = 2.09250061595466E-15
+ ua = -3.382231773605618E-11 lua = -4.49606617112804E-16 wua = -1.427866843597578E-15
+ pua = 2.879320908998649E-22 ub = 1.27558924942704E-18 lub = 3.356660937252002E-25
+ wub = 1.274699373759166E-24 pub = -3.029558420751949E-31 uc = 3.911790161968759E-11
+ luc = 2.503039196218389E-18 wuc = 2.951850404707297E-17 puc = -8.462100869580823E-24
+ ud = 0 up = 0 lp = 1
+ eu = 1.67 vsat = 1.671318384275439E5 lvsat = 3.524244940204454E-4
+ wvsat = 0.023578900102848 pvsat = -9.545537308672942E-9 a0 = 2.844339566190761
+ la0 = -3.071471200444923E-7 wa0 = -2.22891918054084E-6 pa0 = 5.09990165783581E-13
+ ags = 2.063474714004 lags = -4.662421116292038E-7 wags = -1.547404333299792E-6
+ pags = 3.49636009109088E-13 b0 = 0 b1 = 0
+ keta = -1.300488037680807E-3 lketa = -7.87184268154302E-9 wketa = 2.44576963758958E-8
+ pketa = -3.59135274511042E-15 a1 = 0 a2 = 0.38689047
+ rdsw = 103.65 rdswmin = 0 rdw = 0
+ rdwmin = 0 rsw = 0 rswmin = 0
+ prwb = 0 prwg = 0 wr = 1
+ voff = -0.101374184680968 lvoff = -2.009826610000286E-9 wvoff = -2.993828514006634E-8
+ pvoff = 6.474256030176412E-15 voffl = 0 minv = 0
+ nfactor = 2.6731578722336 lnfactor = -5.215358324451204E-8 wnfactor = -5.546849917712932E-7
+ pnfactor = 1.545871190720805E-13 eta0 = -0.01212141499873 leta0 = 5.164790220517678E-9
+ weta0 = 1.392423588565413E-8 peta0 = -4.831445976296357E-15 etab = 0.020937960677445
+ letab = -1.000695102376594E-8 wetab = -1.270028456708572E-8 petab = 6.027669514795147E-15
+ dsub = 1.701534850592136 ldsub = -3.33895512139327E-7 wdsub = -1.075846621520488E-7
+ pdsub = 5.120491995126763E-14 cit = 7.142006000000002E-6 lcit = -1.0194877557E-12
+ wcit = -6.314633688E-12 pcit = 3.0054499038036E-18 cdsc = 3.8556E-37
+ cdscb = -1.1484E-4 cdscd = 4.7984E-6 pclm = 0.289001480567192
+ lpclm = -4.475491385955072E-9 wpclm = -1.664473890096981E-7 ppclm = 9.96382741102458E-14
+ pdiblc1 = 0.39 pdiblc2 = 6.502930906079998E-3 lpdiblc2 = 2.905883546371225E-9
+ wpdiblc2 = -3.458943545523839E-9 ppdiblc2 = -7.282806206896889E-16 pdiblcb = 0
+ drout = 3.4946 pscbe1 = 4.5E8 pscbe2 = 1E-8
+ pvag = 0 delta = 0.01 fprout = 0
+ pdits = 1.4427E-15 pditsl = 0 pditsd = 0
+ lambda = 0 vtl = 0 lc = 0
+ xn = 0 alpha0 = -1.890320172961904E-3 lalpha0 = 9.448465369804022E-10
+ walpha0 = 8.332636244961409E-10 palpha0 = -3.758464896329606E-16 alpha1 = 0
+ beta0 = 16.951384118003997 lbeta0 = 3.112142704333397E-6 wbeta0 = 2.112909345233808E-6
+ pbeta0 = -6.472717239825667E-13 aigbacc = 1 bigbacc = 0
+ cigbacc = 0 nigbacc = 1 aigbinv = 0.35
+ bigbinv = 0.03 cigbinv = 6E-3 eigbinv = 1.1
+ nigbinv = 3 aigc = 0.43 bigc = 0.054
+ cigc = 0.075 aigsd = 0.43 bigsd = 0.054
+ cigsd = 0.075 dlcig = 0 nigc = 1
+ poxedge = 1 pigcd = 1 ntox = 1
+ toxref = 4.148E-9 agidl = 0 bgidl = 2.3E9
+ cgidl = 0.5 egidl = 0.8 noia = 9E41
+ noib = 1E27 noic = 8E11 em = 4.1E7
+ af = 1 ef = 1.2 kf = 0
+ lintnoi = -3E-7 tnoia = 2.5E7 tnoib = 9.9E6
+ ntnoi = 1 rnoia = 0.912 rnoib = 0.26
+ xpart = 0 cgso = {2.392894381E-10/sw_func_tox_lv_ratio} cgdo = {2.392894381E-10/sw_func_tox_lv_ratio}
+ cgbo = {1E-14/sw_func_tox_lv_ratio} ckappas = 0.6 cf = 1E-14
+ clc = 1E-7 cle = 0.6 dlc = 1.21071E-8
+ dwc = 2.6E-8 vfbcv = -1 noff = 3.8661
+ voffcv = -0.16994 acde = 0.38008 moin = 23.81
+ cgsl = {2.310725E-11/sw_func_tox_lv_ratio} cgdl = {2.310725E-11/sw_func_tox_lv_ratio} ijthsrev = 0.1
+ ijthsfwd = 0.1 xjbvs = 1 bvs = 11.9
+ jss = 2.75E-3 jsws = 6E-10 cjs = {1.210E-03*sw_func_nsd_pw_cj}
+ mjs = 0.42197 mjsws = 1E-3 cjsws = {3.230311424E-11*sw_func_nsd_pw_cj}
+ cjswgs = {1.795291232E-10*sw_func_nsd_pw_cj} mjswgs = 0.8 pbs = 0.7477
+ pbsws = 0.1 pbswgs = 0.79644 xrcrg1 = 12
+ xrcrg2 = 1 rbpb = 50 rbpd = 50
+ rbps = 50 rbdb = 50 rbsb = 50
+ gbmin = 1E-12 tnom = 30 ute = -1.4923399698
+ lute = -1.1697396030369E-7 wute = 2.507795495304E-7 pute = 1.553817600266461E-13
+ kt1 = -0.235959719504 lkt1 = -7.896048812071173E-9 wkt1 = -3.244358459020787E-8
+ pkt1 = 7.261166967589451E-15 kt1l = 0 kt2 = -0.0233784172444
+ lkt2 = 1.718735049972179E-9 wkt2 = -2.14641083987088E-8 pkt2 = 2.983209574515454E-15
+ ua1 = -2.038502996599996E-11 lua1 = -1.129409312666824E-16 wua1 = 1.680748342887768E-15
+ pua1 = -2.452747666494108E-23 ub1 = 5.293565084632003E-19 lub1 = -6.751402373060063E-27
+ wub1 = -2.097710505151114E-24 pub1 = 1.829633748838325E-31 uc1 = 5.382616253912004E-11
+ luc1 = -2.297768494869417E-17 wuc1 = -7.834513040292578E-17 puc1 = 2.950305908968612E-23
+ at = 7.584699045799999E4 lat = -4.048231018985098E-3 wat = 0.029470269660216
+ pat = -7.684935404025805E-9 prt = 0 njs = 1.2928
+ xtis = 2 tpb = 1.2287E-3 tpbsw = 0
+ tpbswg = 0 tcj = 7.92E-4 tcjsw = 1E-5
+ tcjswg = 0 tvoff = 0 tvfbsdoff = 0
+ saref = 1.74E-6 sbref = 1.74E-6 wlod = 0
+ ku0 = -2.7E-8 kvsat = 0.2 kvth0 = 7.9E-9
+ tku0 = 0 llodku0 = 0 wlodku0 = 1
+ llodvth = 0 wlodvth = 1 lku0 = 0
+ wku0 = 0 pku0 = 0 lkvth0 = 0
+ wkvth0 = 3E-7 pkvth0 = 0 stk2 = 0
+ lodk2 = 1 steta0 = 0 lodeta0 = 1

.model nlowvt_model.31 nmos
+ level = 54 lmin = 1.8E-7 lmax = 2.5E-7 wmin = 1E-6
+ wmax = 3E-6 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 4.148E-9
+ toxm = 4.148E-9 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 9.999999999999999E22 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {2.6E-8+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {1.2025E-8-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = -1.33E-8 dwb = -1.08E-8 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = 0.542583053185872 lvth0 = -4.250118998523668E-8
+ wvth0 = 7.542728030436521E-8 pvth0 = -1.642565536249254E-14 vfb = 0
+ k1 = 0.386836199729457 lk1 = 4.485035607919113E-8 wk1 = -7.157594991495416E-8
+ pk1 = 1.94235045424411E-14 k2 = -0.021684652994014 lk2 = -1.219435935059446E-8
+ wk2 = 2.279724006706273E-8 pk2 = -5.301754070018006E-15 k3 = 1.65
+ k3b = 1.6 w0 = 1E-7 lpe0 = 2.3802E-7
+ lpeb = -4.9152E-8 vbm = -3 dvtp0 = 0
+ dvtp1 = 0 dvt0 = 0.07665 dvt1 = 0.1252
+ dvt2 = -0.05637 dvt0w = 0 dvt1w = 5.3E6
+ dvt2w = -0.032 vfbsdoff = 0 u0 = 0.030463395807799
+ lu0 = -2.056007076911188E-9 wu0 = -4.442513287221621E-9 pu0 = 2.600158011115919E-16
+ ua = -1.545900105424942E-9 lua = -1.079526409845004E-16 wua = -4.433606652608692E-16
+ pua = 6.54829199046855E-23 ub = 2.800141572552628E-18 lub = -8.806503685026326E-27
+ wub = 3.803390492931375E-25 pub = -1.008751267620958E-31 uc = 6.65613067966257E-11
+ luc = -3.697798203510779E-18 wuc = -2.74621462798331E-19 puc = -1.730344160625404E-24
+ ud = 0 up = 0 lp = 1
+ eu = 1.67 vsat = 1.758516808470715E5 lvsat = -1.617823900671804E-3
+ wvsat = -0.049376985328167 pvsat = 6.9388450044649E-9 a0 = 4.793305784804429
+ la0 = -7.475160371402505E-7 wa0 = 9.09410991482587E-8 pa0 = -1.418226441217094E-14
+ ags = -2.59273113 lags = 5.858275988235E-7 wags = 1.463157298114284E-7
+ pags = -3.306003915089223E-14 b0 = 0 b1 = 0
+ keta = 0.139137388560457 lketa = -3.960378089889229E-8 wketa = 2.463304646035197E-9
+ pketa = 1.378280066251582E-15 a1 = 0 a2 = 0.38689047
+ rdsw = 103.65 rdswmin = 0 rdw = 0
+ rdwmin = 0 rsw = 0 rswmin = 0
+ prwb = 0 prwg = 0 wr = 1
+ voff = -0.145363203121357 lvoff = 7.929492106605653E-9 wvoff = -1.794408637568481E-8
+ pvoff = 3.764166819364406E-15 voffl = 0 minv = 0
+ nfactor = 1.407256058361571 lnfactor = 2.33876931599873E-7 wnfactor = -2.26807034055341E-7
+ pnfactor = 8.050309452616112E-14 eta0 = -0.15010169166732 leta0 = 3.634143373378572E-8
+ weta0 = -5.990410890468526E-9 peta0 = -3.317315372314437E-16 etab = -0.047833289392742
+ letab = 5.531912929592695E-9 wetab = 6.121793985604587E-8 petab = -1.067415329361143E-14
+ dsub = -0.021268339815843 ldsub = 5.53718687333557E-8 wdsub = 3.734448208346762E-7
+ pdsub = -5.748369172958285E-14 cit = -2.650021428571428E-6 lcit = 1.193020841785715E-12
+ wcit = 2.255226317142857E-11 pcit = -3.517025441584286E-18 cdsc = 3.8556E-37
+ cdscb = -1.1484E-4 cdscd = 4.7984E-6 pclm = 0.432211022931457
+ lpclm = -3.683368748316073E-8 wpclm = 7.859248129181217E-7 ppclm = -1.155502249153451E-13
+ pdiblc1 = -0.959235848066286 lpdiblc1 = 3.048598398705773E-7 wpdiblc1 = -9.249644604589565E-9
+ ppdiblc1 = 2.089957198407012E-15 pdiblc2 = 0.037275314161429 lpdiblc2 = -4.047136450174788E-9
+ wpdiblc2 = -2.807225172217716E-8 ppdiblc2 = 4.833096361825127E-15 pdiblcb = 0
+ drout = 3.4946 pscbe1 = 4.5E8 pscbe2 = 1E-8
+ pvag = 0 delta = 0.01 fprout = 0
+ pdits = 1.4427E-15 pditsl = 0 pditsd = 0
+ lambda = 0 vtl = 0 lc = 0
+ xn = 0 alpha0 = 6.105770535162385E-3 lalpha0 = -8.61870158520281E-10
+ walpha0 = -2.453489725346055E-9 palpha0 = 3.667954297638836E-16 alpha1 = 0
+ beta0 = 35.02598114939001 lbeta0 = -9.71812494908272E-7 wbeta0 = -1.472413386707443E-6
+ pbeta0 = 1.628319472995589E-13 aigbacc = 1 bigbacc = 0
+ cigbacc = 0 nigbacc = 1 aigbinv = 0.35
+ bigbinv = 0.03 cigbinv = 6E-3 eigbinv = 1.1
+ nigbinv = 3 aigc = 0.43 bigc = 0.054
+ cigc = 0.075 aigsd = 0.43 bigsd = 0.054
+ cigsd = 0.075 dlcig = 0 nigc = 1
+ poxedge = 1 pigcd = 1 ntox = 1
+ toxref = 4.148E-9 agidl = 0 bgidl = 2.3E9
+ cgidl = 0.5 egidl = 0.8 noia = 9E41
+ noib = 1E27 noic = 8E11 em = 4.1E7
+ af = 1 ef = 1.2 kf = 0
+ lintnoi = -3E-7 tnoia = 2.5E7 tnoib = 9.9E6
+ ntnoi = 1 rnoia = 0.912 rnoib = 0.26
+ xpart = 0 cgso = {2.392894381E-10/sw_func_tox_lv_ratio} cgdo = {2.392894381E-10/sw_func_tox_lv_ratio}
+ cgbo = {1E-14/sw_func_tox_lv_ratio} ckappas = 0.6 cf = 1E-14
+ clc = 1E-7 cle = 0.6 dlc = 1.21071E-8
+ dwc = 2.6E-8 vfbcv = -1 noff = 3.8661
+ voffcv = -0.16994 acde = 0.38008 moin = 23.81
+ cgsl = {2.310725E-11/sw_func_tox_lv_ratio} cgdl = {2.310725E-11/sw_func_tox_lv_ratio} ijthsrev = 0.1
+ ijthsfwd = 0.1 xjbvs = 1 bvs = 11.9
+ jss = 2.75E-3 jsws = 6E-10 cjs = {1.210E-03*sw_func_nsd_pw_cj}
+ mjs = 0.42197 mjsws = 1E-3 cjsws = {3.230311424E-11*sw_func_nsd_pw_cj}
+ cjswgs = {1.795291232E-10*sw_func_nsd_pw_cj} mjswgs = 0.8 pbs = 0.7477
+ pbsws = 0.1 pbswgs = 0.79644 xrcrg1 = 12
+ xrcrg2 = 1 rbpb = 50 rbpd = 50
+ rbps = 50 rbdb = 50 rbsb = 50
+ gbmin = 1E-12 tnom = 30 ute = -2.685764403142858
+ lute = 1.526802904101286E-7 wute = 3.140668991893715E-6 pute = -4.975887594753447E-13
+ kt1 = -0.202390780671428 lkt1 = -1.548095054129075E-8 wkt1 = 4.33110250508544E-9
+ pkt1 = -1.048073581592072E-15 kt1l = 0 kt2 = -1.225288610000003E-3
+ lkt2 = -3.286764364970499E-9 wkt2 = -2.971352149486285E-8 pkt2 = 4.847164463591461E-15
+ ua1 = -1.849359817118572E-9 lua1 = 3.003159218904413E-16 wua1 = 5.739893387256977E-15
+ pua1 = -9.41691299440164E-22 ub1 = 1.322003066517142E-18 lub1 = -1.858498921653485E-25
+ wub1 = -4.817760507915394E-24 pub1 = 7.975586730084217E-31 uc1 = -1.235954070271429E-10
+ luc1 = 1.711071869480293E-17 wuc1 = 1.1670992020116E-16 puc1 = -1.456962959430706E-23
+ at = 3.384537703714286E4 lat = 5.44203353345757E-3 wat = -0.025841228539783
+ pat = 4.812697614263937E-9 prt = 0 njs = 1.2928
+ xtis = 2 tpb = 1.2287E-3 tpbsw = 0
+ tpbswg = 0 tcj = 7.92E-4 tcjsw = 1E-5
+ tcjswg = 0 tvoff = 0 tvfbsdoff = 0
+ saref = 1.25E-6 sbref = 1.24E-6 wlod = 0
+ ku0 = -2.7E-8 kvsat = 0.2 kvth0 = 7.9E-9
+ tku0 = 0 llodku0 = 0 wlodku0 = 1
+ llodvth = 0 wlodvth = 1 lku0 = 0
+ wku0 = 0 pku0 = 0 lkvth0 = 0
+ wkvth0 = 3E-7 pkvth0 = 0 stk2 = 0
+ lodk2 = 1 steta0 = 0 lodeta0 = 1

.model nlowvt_model.32 nmos
+ level = 54 lmin = 1.5E-7 lmax = 1.8E-7 wmin = 1E-6
+ wmax = 3E-6 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 4.148E-9
+ toxm = 4.148E-9 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 9.999999999999999E22 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {2.6E-8+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {1.2025E-8-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = -1.33E-8 dwb = -1.08E-8 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = 0.478426385228733 lvth0 = -3.249595761732098E-8
+ wvth0 = -3.521460050676393E-7 pvth0 = 5.025439849127156E-14 vfb = 0
+ k1 = 0.813026207933334 lk1 = -2.161397570020336E-8 wk1 = 1.910721890792E-7
+ pk1 = -2.153647273369724E-14 k2 = -0.1729664809168 lk2 = 1.139804171396395E-8
+ wk2 = -3.522172340145369E-8 pk2 = 3.746303282897128E-15 k3 = 1.65
+ k3b = 1.6 w0 = 1E-7 lpe0 = 2.3802E-7
+ lpeb = -4.9152E-8 vbm = -3 dvtp0 = 0
+ dvtp1 = 0 dvt0 = 0.07665 dvt1 = 0.1252
+ dvt2 = -0.05637 dvt0w = 0 dvt1w = 5.3E6
+ dvt2w = -0.032 vfbsdoff = 0 u0 = 0.039556021068067
+ lu0 = -3.474001986249996E-9 wu0 = -3.466072868032719E-8 pu0 = 4.972546491666406E-15
+ ua = -1.116456654239469E-9 lua = -1.749243471968749E-16 wua = -1.700256905231385E-15
+ pua = 2.614958885280874E-22 ub = 2.9728711821452E-18 lub = -3.574368630098797E-26
+ wub = -2.904774718440497E-25 pub = 3.738709709248492E-33 uc = 6.99307146511197E-11
+ luc = -4.223257358419115E-18 wuc = 4.730566137205255E-17 puc = -9.150489268720398E-24
+ ud = 0 up = 0 lp = 1
+ eu = 1.67 vsat = 1.472347834944E5 lvsat = 2.844981241477322E-3
+ wvsat = 0.019184922485309 pvsat = -3.753384519046597E-9 a0 = 0
+ ags = 0.809520953999999 lags = 5.524638632370011E-8 wags = -3.320168903919992E-7
+ pags = 4.153593296983229E-14 b0 = 0 b1 = 0
+ keta = 0.4917868334665 lketa = -9.459946183198973E-8 wketa = -9.732738134308423E-7
+ pketa = 1.535444836303406E-13 a1 = 0 a2 = 0.38689047
+ rdsw = 103.65 rdswmin = 0 rdw = 0
+ rdwmin = 0 rsw = 0 rswmin = 0
+ prwb = 0 prwg = 0 wr = 1
+ voff = -0.206349480152747 lvoff = 1.744030200965084E-8 wvoff = 2.114494578476438E-7
+ pvoff = -3.20097564022637E-14 voffl = 0 minv = 0
+ nfactor = 0.243577716870001 lnfactor = 4.153525689554833E-7 wnfactor = 2.261990092701238E-6
+ pnfactor = -3.076248173915273E-13 eta0 = 0.036916430463633 leta0 = 7.175957587463482E-9
+ weta0 = 1.403810407933956E-7 peta0 = -2.315835942733005E-14 etab = -0.08750958174033
+ letab = 1.171943072119906E-8 wetab = 3.097686623667283E-8 petab = -5.958057862670209E-15
+ dsub = 0.6436023713025 ldsub = -4.831471866554986E-8 wdsub = 2.516760265283012E-8
+ pdsub = -3.169859554123953E-15 cit = -1.599166666666667E-5 lcit = 3.273650416666667E-12
+ cdsc = 3.8556E-37 cdscb = -1.1484E-4 cdscd = 4.7984E-6
+ pclm = 0.636703524933334 lpclm = -6.872429317035338E-8 wpclm = -7.186093194368002E-7
+ ppclm = 1.19081873025405E-13 pdiblc1 = 0.8776942606926 lpdiblc1 = 1.839058940962898E-8
+ wpdiblc1 = 3.150246104542147E-7 ppdiblc1 = -4.848061287801351E-14 pdiblc2 = 0.03776610966
+ lpdiblc2 = -4.123676008177001E-9 wpdiblc2 = 5.171823328319991E-9 ppdiblc2 = -3.51317142299903E-16
+ pdiblcb = 0 drout = 3.4946 pscbe1 = 4.5E8
+ pscbe2 = 1E-8 pvag = 0 delta = 0.01
+ fprout = 0 pdits = 1.4427E-15 pditsl = 0
+ pditsd = 0 lambda = 0 vtl = 0
+ lc = 0 xn = 0 alpha0 = 1.311563822895433E-3
+ lalpha0 = -1.142136217422498E-10 walpha0 = 3.439216820155293E-10 palpha0 = -6.946087921415555E-17
+ alpha1 = 0 beta0 = 30.139633958063335 lbeta0 = -2.097866504208765E-7
+ wbeta0 = 4.093810540075963E-6 pbeta0 = -7.052206740823133E-13 aigbacc = 1
+ bigbacc = 0 cigbacc = 0 nigbacc = 1
+ aigbinv = 0.35 bigbinv = 0.03 cigbinv = 6E-3
+ eigbinv = 1.1 nigbinv = 3 aigc = 0.43
+ bigc = 0.054 cigc = 0.075 aigsd = 0.43
+ bigsd = 0.054 cigsd = 0.075 dlcig = 0
+ nigc = 1 poxedge = 1 pigcd = 1
+ ntox = 1 toxref = 4.148E-9 agidl = 0
+ bgidl = 2.3E9 cgidl = 0.5 egidl = 0.8
+ noia = 9E41 noib = 1E27 noic = 8E11
+ em = 4.1E7 af = 1 ef = 1.2
+ kf = 0 lintnoi = -3E-7 tnoia = 2.5E7
+ tnoib = 9.9E6 ntnoi = 1 rnoia = 0.912
+ rnoib = 0.26 xpart = 0 cgso = {2.392894381E-10/sw_func_tox_lv_ratio}
+ cgdo = {2.392894381E-10/sw_func_tox_lv_ratio} cgbo = {1E-14/sw_func_tox_lv_ratio} ckappas = 0.6
+ cf = 1E-14 clc = 1E-7 cle = 0.6
+ dlc = 1.21071E-8 dwc = 2.6E-8 vfbcv = -1
+ noff = 3.8661 voffcv = -0.16994 acde = 0.38008
+ moin = 23.81 cgsl = {2.310725E-11/sw_func_tox_lv_ratio} cgdl = {2.310725E-11/sw_func_tox_lv_ratio}
+ ijthsrev = 0.1 ijthsfwd = 0.1 xjbvs = 1
+ bvs = 11.9 jss = 2.75E-3 jsws = 6E-10
+ cjs = {1.210E-03*sw_func_nsd_pw_cj} mjs = 0.42197 mjsws = 1E-3
+ cjsws = {3.230311424E-11*sw_func_nsd_pw_cj} cjswgs = {1.795291232E-10*sw_func_nsd_pw_cj} mjswgs = 0.8
+ pbs = 0.7477 pbsws = 0.1 pbswgs = 0.79644
+ xrcrg1 = 12 xrcrg2 = 1 rbpb = 50
+ rbpd = 50 rbps = 50 rbdb = 50
+ rbsb = 50 gbmin = 1E-12 tnom = 30
+ ute = -1.870538851 lute = 2.554586555345002E-8 wute = -3.134332732519998E-7
+ pute = 4.107848877412934E-14 kt1 = 0.050186567133333 lkt1 = -5.487038793144334E-8
+ wkt1 = -3.800779274424E-7 pkt1 = 5.890051463871827E-14 kt1l = 0
+ kt2 = -0.059604701205667 lkt2 = 5.817505029323716E-9 wkt2 = -1.474212391902801E-8
+ pkt2 = 2.512375011640018E-15 ua1 = -7.706839094400003E-10 lua1 = 1.32096414087968E-16
+ wua1 = -3.179124850879761E-18 pua1 = -4.60591411769437E-23 ub1 = 1.915012120083333E-18
+ lub1 = -2.783296540689957E-25 wub1 = -1.124297367039E-24 pub1 = 2.21563096188748E-31
+ uc1 = 1.44414679964E-10 luc1 = -2.46854543714658E-17 wuc1 = -3.207419272587202E-17
+ puc1 = 8.63325281666358E-24 at = -3.474074855666667E4 lat = 0.016138039819812
+ wat = 0.10409944255172 pat = -1.545155004245593E-8 prt = 0
+ njs = 1.2928 xtis = 2 tpb = 1.2287E-3
+ tpbsw = 0 tpbswg = 0 tcj = 7.92E-4
+ tcjsw = 1E-5 tcjswg = 0 tvoff = 0
+ tvfbsdoff = 0 saref = 1.1E-6 sbref = 1.1E-6
+ wlod = 0 ku0 = -2.7E-8 kvsat = 0.2
+ kvth0 = 7.9E-9 tku0 = 0 llodku0 = 0
+ wlodku0 = 1 llodvth = 0 wlodvth = 1
+ lku0 = 0 wku0 = 0 pku0 = 0
+ lkvth0 = 0 wkvth0 = 3E-7 pkvth0 = 0
+ stk2 = 0 lodk2 = 1 steta0 = 0
+ lodeta0 = 1

.model nlowvt_model.33 nmos
+ level = 54 lmin = 8E-6 lmax = 2.02E-5 wmin = 4.2E-7
+ wmax = 1E-6 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 4.148E-9
+ toxm = 4.148E-9 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 9.999999999999999E22 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {2.6E-8+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {1.2025E-8-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = -1.33E-8 dwb = -1.08E-8 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = 0.4229525 vfb = 0
+ k1 = 0.53326 k2 = -0.057410608 k3 = 1.65
+ k3b = 1.6 w0 = 1E-7 lpe0 = 2.3802E-7
+ lpeb = -4.9152E-8 vbm = -3 dvtp0 = 0
+ dvtp1 = 0 dvt0 = 0.07665 dvt1 = 0.1252
+ dvt2 = -0.05637 dvt0w = 0 dvt1w = 5.3E6
+ dvt2w = -0.032 vfbsdoff = 0 u0 = 0.0312064
+ ua = -9.7927443E-10 ub = 2.30409E-18 uc = 2.2350587E-11
+ ud = 0 up = 0 lp = 1
+ eu = 1.67 vsat = 2.0055E5 a0 = 1.9208155
+ ags = 0.537176 b0 = 0 b1 = 0
+ keta = 0 a1 = 0 a2 = 0.38689047
+ rdsw = 103.65 rdswmin = 0 rdw = 0
+ rdwmin = 0 rsw = 0 rswmin = 0
+ prwb = 0 prwg = 0 wr = 1
+ voff = -0.11023409 voffl = 0 minv = 0
+ nfactor = 1.6893098 eta0 = 0.08 etab = -0.07
+ dsub = 0.56 cit = 1E-5 cdsc = 3.8556E-37
+ cdscb = -1.1484E-4 cdscd = 4.7984E-6 pclm = 0.2
+ pdiblc1 = 0.39 pdiblc2 = 7.5691E-3 pdiblcb = 0
+ drout = 3.4946 pscbe1 = 4.5E8 pscbe2 = 1E-8
+ pvag = 0 delta = 0.01 fprout = 0
+ pdits = 1.4427E-15 pditsl = 0 pditsd = 0
+ lambda = 0 vtl = 0 lc = 0
+ xn = 0 alpha0 = 4.1734937E-5 alpha1 = 0
+ beta0 = 17.793363 aigbacc = 1 bigbacc = 0
+ cigbacc = 0 nigbacc = 1 aigbinv = 0.35
+ bigbinv = 0.03 cigbinv = 6E-3 eigbinv = 1.1
+ nigbinv = 3 aigc = 0.43 bigc = 0.054
+ cigc = 0.075 aigsd = 0.43 bigsd = 0.054
+ cigsd = 0.075 dlcig = 0 nigc = 1
+ poxedge = 1 pigcd = 1 ntox = 1
+ toxref = 4.148E-9 agidl = 0 bgidl = 2.3E9
+ cgidl = 0.5 egidl = 0.8 noia = 9E41
+ noib = 1E27 noic = 8E11 em = 4.1E7
+ af = 1 ef = 1.2 kf = 0
+ lintnoi = -3E-7 tnoia = 2.5E7 tnoib = 9.9E6
+ ntnoi = 1 rnoia = 0.912 rnoib = 0.26
+ xpart = 0 cgso = {2.392894381E-10/sw_func_tox_lv_ratio} cgdo = {2.392894381E-10/sw_func_tox_lv_ratio}
+ cgbo = {1E-14/sw_func_tox_lv_ratio} ckappas = 0.6 cf = 1E-14
+ clc = 1E-7 cle = 0.6 dlc = 1.21071E-8
+ dwc = 2.6E-8 vfbcv = -1 noff = 3.8661
+ voffcv = -0.16994 acde = 0.38008 moin = 23.81
+ cgsl = {2.310725E-11/sw_func_tox_lv_ratio} cgdl = {2.310725E-11/sw_func_tox_lv_ratio} ijthsrev = 0.1
+ ijthsfwd = 0.1 xjbvs = 1 bvs = 11.9
+ jss = 2.75E-3 jsws = 6E-10 cjs = {1.210E-03*sw_func_nsd_pw_cj}
+ mjs = 0.42197 mjsws = 1E-3 cjsws = {3.230311424E-11*sw_func_nsd_pw_cj}
+ cjswgs = {1.795291232E-10*sw_func_nsd_pw_cj} mjswgs = 0.8 pbs = 0.7477
+ pbsws = 0.1 pbswgs = 0.79644 xrcrg1 = 12
+ xrcrg2 = 1 rbpb = 50 rbpd = 50
+ rbps = 50 rbdb = 50 rbsb = 50
+ gbmin = 1E-12 tnom = 30 ute = -1.1808
+ kt1 = -0.25763 kt1l = 0 kt2 = -0.036364
+ ua1 = 1.9636E-9 ub1 = -1.466E-18 uc1 = 6.3418E-11
+ at = 5.823E4 prt = 0 njs = 1.2928
+ xtis = 2 tpb = 1.2287E-3 tpbsw = 0
+ tpbswg = 0 tcj = 7.92E-4 tcjsw = 1E-5
+ tcjswg = 0 tvoff = 0 tvfbsdoff = 0
+ saref = 3E-6 sbref = 3E-6 wlod = 0
+ ku0 = -2.7E-8 kvsat = 0.2 kvth0 = 7.9E-9
+ tku0 = 0 llodku0 = 0 wlodku0 = 1
+ llodvth = 0 wlodvth = 1 lku0 = 0
+ wku0 = 0 pku0 = 0 lkvth0 = 0
+ wkvth0 = 3E-7 pkvth0 = 0 stk2 = 0
+ lodk2 = 1 steta0 = 0 lodeta0 = 1

.model nlowvt_model.34 nmos
+ level = 54 lmin = 4E-6 lmax = 8E-6 wmin = 4.2E-7
+ wmax = 1E-6 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 4.148E-9
+ toxm = 4.148E-9 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 9.999999999999999E22 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {2.6E-8+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {1.2025E-8-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = -1.33E-8 dwb = -1.08E-8 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = 0.4229525 vfb = 0
+ k1 = 0.53326 k2 = -0.057410608 k3 = 1.65
+ k3b = 1.6 w0 = 1E-7 lpe0 = 2.3802E-7
+ lpeb = -4.9152E-8 vbm = -3 dvtp0 = 0
+ dvtp1 = 0 dvt0 = 0.07665 dvt1 = 0.1252
+ dvt2 = -0.05637 dvt0w = 0 dvt1w = 5.3E6
+ dvt2w = -0.032 vfbsdoff = 0 u0 = 0.0312064
+ ua = -9.7927443E-10 ub = 2.30409E-18 uc = 2.2350587E-11
+ ud = 0 up = 0 lp = 1
+ eu = 1.67 vsat = 2.0055E5 a0 = 1.9208155
+ ags = 0.537176 b0 = 0 b1 = 0
+ keta = 0 a1 = 0 a2 = 0.38689047
+ rdsw = 103.65 rdswmin = 0 rdw = 0
+ rdwmin = 0 rsw = 0 rswmin = 0
+ prwb = 0 prwg = 0 wr = 1
+ voff = -0.11023409 voffl = 0 minv = 0
+ nfactor = 1.6893098 eta0 = 0.08 etab = -0.07
+ dsub = 0.56 cit = 1E-5 cdsc = 3.8556E-37
+ cdscb = -1.1484E-4 cdscd = 4.7984E-6 pclm = 0.2
+ pdiblc1 = 0.39 pdiblc2 = 7.5691E-3 pdiblcb = 0
+ drout = 3.4946 pscbe1 = 4.5E8 pscbe2 = 1E-8
+ pvag = 0 delta = 0.01 fprout = 0
+ pdits = 1.4427E-15 pditsl = 0 pditsd = 0
+ lambda = 0 vtl = 0 lc = 0
+ xn = 0 alpha0 = 4.1734937E-5 alpha1 = 0
+ beta0 = 17.793363 aigbacc = 1 bigbacc = 0
+ cigbacc = 0 nigbacc = 1 aigbinv = 0.35
+ bigbinv = 0.03 cigbinv = 6E-3 eigbinv = 1.1
+ nigbinv = 3 aigc = 0.43 bigc = 0.054
+ cigc = 0.075 aigsd = 0.43 bigsd = 0.054
+ cigsd = 0.075 dlcig = 0 nigc = 1
+ poxedge = 1 pigcd = 1 ntox = 1
+ toxref = 4.148E-9 agidl = 0 bgidl = 2.3E9
+ cgidl = 0.5 egidl = 0.8 noia = 9E41
+ noib = 1E27 noic = 8E11 em = 4.1E7
+ af = 1 ef = 1.2 kf = 0
+ lintnoi = -3E-7 tnoia = 2.5E7 tnoib = 9.9E6
+ ntnoi = 1 rnoia = 0.912 rnoib = 0.26
+ xpart = 0 cgso = {2.392894381E-10/sw_func_tox_lv_ratio} cgdo = {2.392894381E-10/sw_func_tox_lv_ratio}
+ cgbo = {1E-14/sw_func_tox_lv_ratio} ckappas = 0.6 cf = 1E-14
+ clc = 1E-7 cle = 0.6 dlc = 1.21071E-8
+ dwc = 2.6E-8 vfbcv = -1 noff = 3.8661
+ voffcv = -0.16994 acde = 0.38008 moin = 23.81
+ cgsl = {2.310725E-11/sw_func_tox_lv_ratio} cgdl = {2.310725E-11/sw_func_tox_lv_ratio} ijthsrev = 0.1
+ ijthsfwd = 0.1 xjbvs = 1 bvs = 11.9
+ jss = 2.75E-3 jsws = 6E-10 cjs = {1.210E-03*sw_func_nsd_pw_cj}
+ mjs = 0.42197 mjsws = 1E-3 cjsws = {3.230311424E-11*sw_func_nsd_pw_cj}
+ cjswgs = {1.795291232E-10*sw_func_nsd_pw_cj} mjswgs = 0.8 pbs = 0.7477
+ pbsws = 0.1 pbswgs = 0.79644 xrcrg1 = 12
+ xrcrg2 = 1 rbpb = 50 rbpd = 50
+ rbps = 50 rbdb = 50 rbsb = 50
+ gbmin = 1E-12 tnom = 30 ute = -1.1808
+ kt1 = -0.25763 kt1l = 0 kt2 = -0.036364
+ ua1 = 1.9636E-9 ub1 = -1.466E-18 uc1 = 6.3418E-11
+ at = 5.823E4 prt = 0 njs = 1.2928
+ xtis = 2 tpb = 1.2287E-3 tpbsw = 0
+ tpbswg = 0 tcj = 7.92E-4 tcjsw = 1E-5
+ tcjswg = 0 tvoff = 0 tvfbsdoff = 0
+ saref = 3E-6 sbref = 3E-6 wlod = 0
+ ku0 = -2.7E-8 kvsat = 0.2 kvth0 = 7.9E-9
+ tku0 = 0 llodku0 = 0 wlodku0 = 1
+ llodvth = 0 wlodvth = 1 lku0 = 0
+ wku0 = 0 pku0 = 0 lkvth0 = 0
+ wkvth0 = 3E-7 pkvth0 = 0 stk2 = 0
+ lodk2 = 1 steta0 = 0 lodeta0 = 1

.model nlowvt_model.35 nmos
+ level = 54 lmin = 2E-6 lmax = 4E-6 wmin = 4.2E-7
+ wmax = 1E-6 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 4.148E-9
+ toxm = 4.148E-9 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 9.999999999999999E22 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {2.6E-8+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {1.2025E-8-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = -1.33E-8 dwb = -1.08E-8 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = 0.40400458327373 lvth0 = 7.533596950781147E-8
+ wvth0 = 7.66123933689357E-9 pvth0 = -3.046070454152199E-14 vfb = 0
+ k1 = 0.643847734324712 lk1 = -4.396913022883408E-7 wk1 = -3.428307154082757E-8
+ pk1 = 1.363077782927534E-13 k2 = -0.102202454835322 lk2 = 1.780901434248973E-7
+ wk2 = 1.476467629521256E-8 pk2 = -5.870361471595039E-14 k3 = 1.65
+ k3b = 1.6 w0 = 1E-7 lpe0 = 2.3802E-7
+ lpeb = -4.9152E-8 vbm = -3 dvtp0 = 0
+ dvtp1 = 0 dvt0 = 0.07665 dvt1 = 0.1252
+ dvt2 = -0.05637 dvt0w = 0 dvt1w = 5.3E6
+ dvt2w = -0.032 vfbsdoff = 0 u0 = 0.030704042934416
+ lu0 = 1.997346574908378E-9 wu0 = 2.634014460015539E-10 pu0 = -1.047270979229878E-15
+ ua = -8.119869376501484E-10 lua = -6.65126705208392E-16 wua = -3.694779420322816E-17
+ pua = 1.46902582362325E-22 ub = 2.07591511092816E-18 lub = 9.072119502051797E-25
+ wub = 5.228298430110338E-26 pub = -2.07874531431972E-31 uc = -2.407790188367066E-11
+ luc = 1.845973503770303E-16 wuc = 1.674563951159587E-17 puc = -6.657982541612959E-23
+ ud = 0 up = 0 lp = 1
+ eu = 1.67 vsat = 4.329783050990807E5 lvsat = -0.92412331965869
+ wvsat = -0.072497802678328 pvsat = 2.882476385588999E-7 a0 = 1.957496949687155
+ la0 = -1.458436098836443E-7 wa0 = 2.972075065472698E-8 pa0 = -1.181682185656617E-13
+ ags = -0.687184137994368 lags = 4.867994690658708E-6 wags = 3.043279121184608E-7
+ pags = -1.209992562187394E-12 b0 = 1.663832764735631E-8 lb0 = -6.615315880950633E-14
+ wb0 = -1.577313460969378E-14 pb0 = 6.271319455141199E-20 b1 = 4.586588081379302E-10
+ lb1 = -1.823604488216005E-15 wb1 = -4.348085501147581E-16 pb1 = 1.728777054828772E-21
+ keta = 0.265822281095977 lketa = -1.056896098523549E-6 wketa = -8.225945010998589E-8
+ pketa = 3.270594606647984E-13 a1 = 0 a2 = 0.38689047
+ rdsw = 103.65 rdswmin = 0 rdw = 0
+ rdwmin = 0 rsw = 0 rswmin = 0
+ prwb = 0 prwg = 0 wr = 1
+ voff = -0.103356304183205 lvoff = -2.734573251828798E-8 wvoff = -1.45939024618115E-10
+ pvoff = 5.802462649303944E-16 voffl = 0 minv = 0
+ nfactor = 2.22282600341487 lnfactor = -2.121233748967355E-6 wnfactor = -1.647500453470084E-7
+ pnfactor = 6.550379427974379E-13 eta0 = 0.191879449585368 leta0 = -4.448270975789454E-7
+ weta0 = -3.160199435692921E-8 peta0 = 1.256479494634327E-13 etab = -0.167782006063218
+ letab = 3.887763670070519E-7 wetab = 2.760362089793072E-8 petab = -1.097506165091276E-13
+ dsub = 0.752827963101855 ldsub = -7.666743398948213E-7 wdsub = -3.504573042148265E-8
+ pdsub = 1.393400718692939E-13 cit = 1E-5 cdsc = 3.8556E-37
+ cdscb = -1.1484E-4 cdscd = 4.7984E-6 pclm = 0.153379723684482
+ lpclm = 1.853598876166818E-7 wpclm = 1.185521358811061E-8 ppclm = -4.713573646564838E-14
+ pdiblc1 = 0.39 pdiblc2 = 1.629167205534479E-3 lpdiblc2 = 2.361687579415518E-8
+ wpdiblc2 = 1.717097295483312E-9 ppdiblc2 = -6.827092991976874E-15 pdiblcb = 0
+ drout = 3.4946 pscbe1 = 4.5E8 pscbe2 = 1E-8
+ pvag = 0 delta = 0.01 fprout = 0
+ pdits = 1.4427E-15 pditsl = 0 pditsd = 0
+ lambda = 0 vtl = 0 lc = 0
+ xn = 0 alpha0 = -8.217749125803262E-5 lalpha0 = 4.926696191325248E-10
+ walpha0 = 4.001219056483201E-11 palpha0 = -1.590864690762438E-16 alpha1 = 0
+ beta0 = 13.154233423395402 lbeta0 = 1.844494724010105E-5 wbeta0 = 1.215446904059558E-6
+ pbeta0 = -4.832556118195598E-12 aigbacc = 1 bigbacc = 0
+ cigbacc = 0 nigbacc = 1 aigbinv = 0.35
+ bigbinv = 0.03 cigbinv = 6E-3 eigbinv = 1.1
+ nigbinv = 3 aigc = 0.43 bigc = 0.054
+ cigc = 0.075 aigsd = 0.43 bigsd = 0.054
+ cigsd = 0.075 dlcig = 0 nigc = 1
+ poxedge = 1 pigcd = 1 ntox = 1
+ toxref = 4.148E-9 agidl = 0 bgidl = 2.3E9
+ cgidl = 0.5 egidl = 0.8 noia = 9E41
+ noib = 1E27 noic = 8E11 em = 4.1E7
+ af = 1 ef = 1.2 kf = 0
+ lintnoi = -3E-7 tnoia = 2.5E7 tnoib = 9.9E6
+ ntnoi = 1 rnoia = 0.912 rnoib = 0.26
+ xpart = 0 cgso = {2.392894381E-10/sw_func_tox_lv_ratio} cgdo = {2.392894381E-10/sw_func_tox_lv_ratio}
+ cgbo = {1E-14/sw_func_tox_lv_ratio} ckappas = 0.6 cf = 1E-14
+ clc = 1E-7 cle = 0.6 dlc = 1.21071E-8
+ dwc = 2.6E-8 vfbcv = -1 noff = 3.8661
+ voffcv = -0.16994 acde = 0.38008 moin = 23.81
+ cgsl = {2.310725E-11/sw_func_tox_lv_ratio} cgdl = {2.310725E-11/sw_func_tox_lv_ratio} ijthsrev = 0.1
+ ijthsfwd = 0.1 xjbvs = 1 bvs = 11.9
+ jss = 2.75E-3 jsws = 6E-10 cjs = {1.210E-03*sw_func_nsd_pw_cj}
+ mjs = 0.42197 mjsws = 1E-3 cjsws = {3.230311424E-11*sw_func_nsd_pw_cj}
+ cjswgs = {1.795291232E-10*sw_func_nsd_pw_cj} mjswgs = 0.8 pbs = 0.7477
+ pbsws = 0.1 pbswgs = 0.79644 xrcrg1 = 12
+ xrcrg2 = 1 rbpb = 50 rbpd = 50
+ rbps = 50 rbdb = 50 rbsb = 50
+ gbmin = 1E-12 tnom = 30 ute = -1.253788864798851
+ lute = 2.902000769969908E-7 wute = 1.196716549931038E-8 pute = -4.758085166698312E-14
+ kt1 = -0.239613129617816 lkt1 = -7.163417579604447E-8 wkt1 = -6.88041585531047E-9
+ pkt1 = 2.735618941992166E-14 kt1l = 0 kt2 = -0.034241296777184
+ lkt2 = -8.439761878756905E-9 wkt2 = -1.33328743772996E-9 pkt2 = 5.301084188042433E-15
+ ua1 = 1.859859004488506E-9 lua1 = 4.124690111039264E-16 wua1 = 2.0889618934897E-17
+ pua1 = -8.305608040420373E-23 ub1 = -8.632276881206892E-19 lub1 = -2.396592573416545E-24
+ wub1 = -1.702822431715863E-25 pub1 = 6.770336847380686E-31 uc1 = 1.753860372198218E-10
+ luc1 = -4.451793175841506E-16 wuc1 = -3.81409310419611E-17 puc1 = 1.516464347762852E-22
+ at = 7.8391319326092E4 lat = -0.080160397574575 wat = -0.010629205203735
+ pat = 4.226118842979099E-8 prt = 0 njs = 1.2928
+ xtis = 2 tpb = 1.2287E-3 tpbsw = 0
+ tpbswg = 0 tcj = 7.92E-4 tcjsw = 1E-5
+ tcjswg = 0 tvoff = 0 tvfbsdoff = 0
+ saref = 3E-6 sbref = 3E-6 wlod = 0
+ ku0 = -2.7E-8 kvsat = 0.2 kvth0 = 7.9E-9
+ tku0 = 0 llodku0 = 0 wlodku0 = 1
+ llodvth = 0 wlodvth = 1 lku0 = 0
+ wku0 = 0 pku0 = 0 lkvth0 = 0
+ wkvth0 = 3E-7 pkvth0 = 0 stk2 = 0
+ lodk2 = 1 steta0 = 0 lodeta0 = 1

.model nlowvt_model.36 nmos
+ level = 54 lmin = 1E-6 lmax = 2E-6 wmin = 4.2E-7
+ wmax = 1E-6 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 4.148E-9
+ toxm = 4.148E-9 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 9.999999999999999E22 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {2.6E-8+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {1.2025E-8-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = -1.33E-8 dwb = -1.08E-8 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = 0.432261574697298 lvth0 = 1.950156730441362E-8
+ wvth0 = -2.737333506978321E-9 pvth0 = -9.913644530673325E-15 vfb = 0
+ k1 = 0.399794975136782 lk1 = 4.254474722905108E-8 wk1 = 5.552834384033103E-8
+ pk1 = -4.115508792964693E-14 k2 = 1.407966400491657E-3 lk2 = -2.66388684160081E-8
+ wk2 = -2.336395871956609E-8 pk2 = 1.663666164150149E-14 k3 = 1.65
+ k3b = 1.6 w0 = 1E-7 lpe0 = 2.3802E-7
+ lpeb = -4.9152E-8 vbm = -3 dvtp0 = 0
+ dvtp1 = 0 dvt0 = 0.07665 dvt1 = 0.1252
+ dvt2 = -0.05637 dvt0w = 0 dvt1w = 5.3E6
+ dvt2w = -0.032 vfbsdoff = 0 u0 = 0.039151637572825
+ lu0 = -1.469467805085586E-8 wu0 = -2.84531338093297E-9 pu0 = 5.095394083051395E-15
+ ua = -5.946337063815512E-10 lua = -1.094605822533577E-15 wua = -1.169337833100715E-16
+ pua = 3.049508975379922E-22 ub = 2.440194506647126E-18 lub = 1.87414078234289E-25
+ wub = -8.177183332347561E-26 pub = 5.701108545331491E-32 uc = 8.158161886343954E-11
+ luc = -2.41805796432221E-17 wuc = -2.213706412334069E-17 puc = 1.025045283132331E-23
+ ud = 0 up = 0 lp = 1
+ eu = 1.67 vsat = -1.459689035119542E5 lvsat = 0.219847417196285
+ wvsat = 0.140554770090533 pvsat = -1.327335926037312E-7 a0 = 2.328177998355518
+ la0 = -8.78290827999895E-7 wa0 = -1.066898752552306E-7 pa0 = 1.513723577011189E-13
+ ags = 1.86143313759908 lags = -1.679456150501674E-7 wags = -6.33563245299928E-7
+ pags = 6.432334703134717E-13 b0 = 1.663832764735635E-8 lb0 = -6.615315880950639E-14
+ wb0 = -1.577313460969382E-14 pb0 = 6.271319455141206E-20 b1 = 4.586588081379321E-10
+ lb1 = -1.823604488216008E-15 wb1 = -4.348085501147597E-16 pb1 = 1.728777054828776E-21
+ keta = -0.432670645802298 lketa = 3.232910003810976E-7 wketa = 1.747859469885786E-7
+ pketa = -1.808493917321102E-13 a1 = 0 a2 = 0.38689047
+ rdsw = 103.65 rdswmin = 0 rdw = 0
+ rdwmin = 0 rsw = 0 rswmin = 0
+ prwb = 0 prwg = 0 wr = 1
+ voff = -0.128484281975363 lvoff = 2.230589520012831E-8 wvoff = 9.10115680289648E-9
+ pvoff = -1.769155273544707E-14 voffl = 0 minv = 0
+ nfactor = 0.072802324138652 lnfactor = 2.127105540098489E-6 wnfactor = 6.264586686266399E-7
+ pnfactor = -9.083509155787926E-13 eta0 = -0.066334653011335 leta0 = 6.539105844701132E-8
+ weta0 = 6.342079539865789E-8 peta0 = -6.211233195411966E-14 etab = 0.058000290428412
+ letab = -5.735816174558451E-8 wetab = -5.548426421098854E-8 petab = 5.442689007184139E-14
+ dsub = -0.031732182622679 ldsub = 7.835772800495728E-7 wdsub = 2.536724032051458E-7
+ pdsub = -4.311525242702426E-13 cit = 1.79758672413793E-5 lcit = -1.575991487560344E-11
+ wcit = -2.935119144827576E-12 pcit = 5.79964867422206E-18 cdsc = 3.8556E-37
+ cdscb = -1.1484E-4 cdscd = 4.7984E-6 pclm = 0.301645299417242
+ lpclm = -1.076054767524641E-7 wpclm = -4.270651828154533E-8 ppclm = 6.067551762219829E-14
+ pdiblc1 = 0.39 pdiblc2 = 0.010509926561862 lpdiblc2 = 6.068939344019674E-9
+ wpdiblc2 = -1.551022147645245E-9 ppdiblc2 = -3.694523783270023E-16 pdiblcb = 0
+ drout = 3.4946 pscbe1 = 4.5E8 pscbe2 = 1E-8
+ pvag = 0 delta = 0.01 fprout = 0
+ pdits = 1.4427E-15 pditsl = 0 pditsd = 0
+ lambda = 0 vtl = 0 lc = 0
+ xn = 0 alpha0 = 3.099688777322006E-4 lalpha0 = -2.821919986737267E-10
+ walpha0 = -1.042976732235738E-10 palpha0 = 1.260626062764568E-16 alpha1 = 0
+ beta0 = 24.8622273032885 lbeta0 = -4.689463266873723E-6 wbeta0 = -3.0930948437411E-6
+ pbeta0 = 3.680906948371112E-12 aigbacc = 1 bigbacc = 0
+ cigbacc = 0 nigbacc = 1 aigbinv = 0.35
+ bigbinv = 0.03 cigbinv = 6E-3 eigbinv = 1.1
+ nigbinv = 3 aigc = 0.43 bigc = 0.054
+ cigc = 0.075 aigsd = 0.43 bigsd = 0.054
+ cigsd = 0.075 dlcig = 0 nigc = 1
+ poxedge = 1 pigcd = 1 ntox = 1
+ toxref = 4.148E-9 agidl = 0 bgidl = 2.3E9
+ cgidl = 0.5 egidl = 0.8 noia = 9E41
+ noib = 1E27 noic = 8E11 em = 4.1E7
+ af = 1 ef = 1.2 kf = 0
+ lintnoi = -3E-7 tnoia = 2.5E7 tnoib = 9.9E6
+ ntnoi = 1 rnoia = 0.912 rnoib = 0.26
+ xpart = 0 cgso = {2.392894381E-10/sw_func_tox_lv_ratio} cgdo = {2.392894381E-10/sw_func_tox_lv_ratio}
+ cgbo = {1E-14/sw_func_tox_lv_ratio} ckappas = 0.6 cf = 1E-14
+ clc = 1E-7 cle = 0.6 dlc = 1.21071E-8
+ dwc = 2.6E-8 vfbcv = -1 noff = 3.8661
+ voffcv = -0.16994 acde = 0.38008 moin = 23.81
+ cgsl = {2.310725E-11/sw_func_tox_lv_ratio} cgdl = {2.310725E-11/sw_func_tox_lv_ratio} ijthsrev = 0.1
+ ijthsfwd = 0.1 xjbvs = 1 bvs = 11.9
+ jss = 2.75E-3 jsws = 6E-10 cjs = {1.210E-03*sw_func_nsd_pw_cj}
+ mjs = 0.42197 mjsws = 1E-3 cjsws = {3.230311424E-11*sw_func_nsd_pw_cj}
+ cjswgs = {1.795291232E-10*sw_func_nsd_pw_cj} mjswgs = 0.8 pbs = 0.7477
+ pbsws = 0.1 pbswgs = 0.79644 xrcrg1 = 12
+ xrcrg2 = 1 rbpb = 50 rbpd = 50
+ rbps = 50 rbdb = 50 rbsb = 50
+ gbmin = 1E-12 tnom = 30 ute = -1.09800661954023
+ lute = -1.761785052178178E-8 wute = -4.536070075586212E-8 pute = 6.5696145659925E-14
+ kt1 = -0.273386999722989 lkt1 = -4.898697161728447E-9 wkt1 = 5.548368343393349E-9
+ pkt1 = 2.797533282492848E-15 kt1l = 0 kt2 = -0.05952766547115
+ lkt2 = 4.152483834208614E-8 wkt2 = 7.972096241650264E-9 pkt2 = -1.308588869322892E-14
+ ua1 = 2.209452306609196E-9 lua1 = -2.783098742214519E-16 wua1 = -1.077607162455182E-16
+ pua1 = 1.711505493955377E-22 ub1 = -2.524013291068964E-18 lub1 = 8.850367387291006E-25
+ wub1 = 4.408868587133791E-25 pub1 = -5.30605902131529E-31 uc1 = 4.490025664149444E-12
+ luc1 = -1.074973435507197E-16 wuc1 = 2.474880121052633E-17 puc1 = 2.737946833198268E-23
+ at = 2.091270453678098E3 lat = 0.070604683994871 wat = 0.017449212781313
+ pat = -1.322036158776534E-8 prt = 0 njs = 1.2928
+ xtis = 2 tpb = 1.2287E-3 tpbsw = 0
+ tpbswg = 0 tcj = 7.92E-4 tcjsw = 1E-5
+ tcjswg = 0 tvoff = 0 tvfbsdoff = 0
+ saref = 3E-6 sbref = 3E-6 wlod = 0
+ ku0 = -2.7E-8 kvsat = 0.2 kvth0 = 7.9E-9
+ tku0 = 0 llodku0 = 0 wlodku0 = 1
+ llodvth = 0 wlodvth = 1 lku0 = 0
+ wku0 = 0 pku0 = 0 lkvth0 = 0
+ wkvth0 = 3E-7 pkvth0 = 0 stk2 = 0
+ lodk2 = 1 steta0 = 0 lodeta0 = 1

.model nlowvt_model.37 nmos
+ level = 54 lmin = 5E-7 lmax = 1E-6 wmin = 4.2E-7
+ wmax = 1E-6 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 4.148E-9
+ toxm = 4.148E-9 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 9.999999999999999E22 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {2.6E-8+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {1.2025E-8-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = -1.33E-8 dwb = -1.08E-8 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = 0.449932663330493 lvth0 = 2.255468352846905E-9
+ wvth0 = -2.881846994987164E-9 pvth0 = -9.772606592051093E-15 vfb = 0
+ k1 = 0.444939542129016 lk1 = -1.514092927020357E-9 wk1 = -2.017648430307378E-9
+ pk1 = 1.500692322688263E-14 k2 = -0.017295236376082 lk2 = -8.385477666211519E-9
+ wk2 = -5.529989784148322E-9 pk2 = -7.684003410194786E-16 k3 = 1.65
+ k3b = 1.6 w0 = 1E-7 lpe0 = 2.3802E-7
+ lpeb = -4.9152E-8 vbm = -3 dvtp0 = 0
+ dvtp1 = 0 dvt0 = 0.07665 dvt1 = 0.1252
+ dvt2 = -0.05637 dvt0w = 0 dvt1w = 5.3E6
+ dvt2w = -0.032 vfbsdoff = 0 u0 = 0.029350328301709
+ lu0 = -5.129090267710535E-9 wu0 = 1.031645363205079E-9 pu0 = 1.311676196709868E-15
+ ua = -1.265948535447975E-9 lua = -4.394361151062008E-16 wua = 7.239210444368393E-17
+ pua = 1.201782973847145E-22 ub = 2.564840245350883E-18 lub = 6.576606954635719E-26
+ wub = -1.371720308637402E-27 pub = -2.145540484351643E-32 uc = 3.55345360065024E-11
+ luc = 2.075907087100571E-17 wuc = -2.503089436929471E-18 puc = -8.911324763879716E-24
+ ud = 0 up = 0 lp = 1
+ eu = 1.67 vsat = -4.846086928127955E4 lvsat = 0.124684451188858
+ wvsat = 0.046710394607413 pvsat = -4.114617435098061E-8 a0 = 2.019812794930463
+ la0 = -5.773418077172128E-7 wa0 = -6.011849136367864E-8 pa0 = 1.059210155921588E-13
+ ags = 3.927687899292514 lags = -2.184506949724874E-6 wags = -7.520449087933039E-7
+ pags = 7.588656497998318E-13 b0 = -6.087193041715727E-8 lb0 = 9.492977548555677E-15
+ wb0 = 5.77065900354651E-14 pb0 = -8.99934271603078E-21 b1 = -1.678020029772917E-9
+ lb1 = 2.616872236430855E-16 wb1 = 1.590762988224725E-15 pb1 = -2.48079488013645E-22
+ keta = -0.26077635826291 lketa = 1.555307704570318E-7 wketa = 3.902734862123869E-8
+ pketa = -4.835578765550479E-14 a1 = 0 a2 = 0.38689047
+ rdsw = 103.65 rdswmin = 0 rdw = 0
+ rdwmin = 0 rsw = 0 rswmin = 0
+ prwb = 0 prwg = 0 wr = 1
+ voff = -0.092731677061406 lvoff = -1.258685956564885E-8 wvoff = -1.432386117985156E-8
+ pvoff = 5.170093564815876E-15 voffl = 0 minv = 0
+ nfactor = 1.80916414705157 lnfactor = 4.325032190266276E-7 wnfactor = -2.358464276329678E-7
+ pnfactor = -6.678425688422848E-14 eta0 = 5.888087402591273E-3 leta0 = -5.094725059960331E-9
+ weta0 = -7.225445949991686E-9 peta0 = 6.834867290094893E-15 etab = -5.100268866479902E-3
+ letab = 4.224829098265197E-9 wetab = 4.074632205130946E-9 petab = -3.699614885470429E-15
+ dsub = 0.113393243502799 ldsub = 6.419421204224119E-7 wdsub = 4.988537460535027E-8
+ pdsub = -2.322665737082722E-13 cit = 1.827586206896549E-6 wcit = 3.00744827586207E-12
+ cdsc = 3.8556E-37 cdscb = -1.1484E-4 cdscd = 4.7984E-6
+ pclm = 0.023758282533389 lpclm = 1.63598357375332E-7 wpclm = 7.646914064234714E-8
+ ppclm = -5.563396670457456E-14 pdiblc1 = 0.347645606391926 lpdiblc1 = 4.13357704418001E-8
+ wpdiblc1 = 4.015196514045443E-8 ppdiblc1 = -3.91863103788265E-14 pdiblc2 = 0.028263509818843
+ lpdiblc2 = -1.125767023563067E-8 wpdiblc2 = -6.234540731382981E-9 ppdiblc2 = 4.20142758347184E-15
+ pdiblcb = 0 drout = 3.4946 pscbe1 = 4.5E8
+ pscbe2 = 1E-8 pvag = 0 delta = 0.01
+ fprout = 0 pdits = 1.4427E-15 pditsl = 0
+ pditsd = 0 lambda = 0 vtl = 0
+ lc = 0 xn = 0 alpha0 = -7.487820553054027E-5
+ lalpha0 = 9.339951223654527E-11 walpha0 = 3.096937032193542E-11 palpha0 = -5.951264871783006E-18
+ alpha1 = 0 beta0 = 15.401708385770327 lbeta0 = 4.543530170678136E-6
+ wbeta0 = 1.923148509292128E-6 pbeta0 = -1.214695752021667E-12 aigbacc = 1
+ bigbacc = 0 cigbacc = 0 nigbacc = 1
+ aigbinv = 0.35 bigbinv = 0.03 cigbinv = 6E-3
+ eigbinv = 1.1 nigbinv = 3 aigc = 0.43
+ bigc = 0.054 cigc = 0.075 aigsd = 0.43
+ bigsd = 0.054 cigsd = 0.075 dlcig = 0
+ nigc = 1 poxedge = 1 pigcd = 1
+ ntox = 1 toxref = 4.148E-9 agidl = 0
+ bgidl = 2.3E9 cgidl = 0.5 egidl = 0.8
+ noia = 9E41 noib = 1E27 noic = 8E11
+ em = 4.1E7 af = 1 ef = 1.2
+ kf = 0 lintnoi = -3E-7 tnoia = 2.5E7
+ tnoib = 9.9E6 ntnoi = 1 rnoia = 0.912
+ rnoib = 0.26 xpart = 0 cgso = {2.392894381E-10/sw_func_tox_lv_ratio}
+ cgdo = {2.392894381E-10/sw_func_tox_lv_ratio} cgbo = {1E-14/sw_func_tox_lv_ratio} ckappas = 0.6
+ cf = 1E-14 clc = 1E-7 cle = 0.6
+ dlc = 1.21071E-8 dwc = 2.6E-8 vfbcv = -1
+ noff = 3.8661 voffcv = -0.16994 acde = 0.38008
+ moin = 23.81 cgsl = {2.310725E-11/sw_func_tox_lv_ratio} cgdl = {2.310725E-11/sw_func_tox_lv_ratio}
+ ijthsrev = 0.1 ijthsfwd = 0.1 xjbvs = 1
+ bvs = 11.9 jss = 2.75E-3 jsws = 6E-10
+ cjs = {1.210E-03*sw_func_nsd_pw_cj} mjs = 0.42197 mjsws = 1E-3
+ cjsws = {3.230311424E-11*sw_func_nsd_pw_cj} cjswgs = {1.795291232E-10*sw_func_nsd_pw_cj} mjswgs = 0.8
+ pbs = 0.7477 pbsws = 0.1 pbswgs = 0.79644
+ xrcrg1 = 12 xrcrg2 = 1 rbpb = 50
+ rbpd = 50 rbps = 50 rbdb = 50
+ rbsb = 50 gbmin = 1E-12 tnom = 30
+ ute = -1.142274387638351 lute = 2.558527775358027E-8 wute = 7.95640830411573E-8
+ pute = -5.62241970867761E-14 kt1 = -0.278248598529016 lkt1 = -1.540198069860482E-10
+ wkt1 = 9.30299278550725E-9 pkt1 = -8.667924417882124E-16 kt1l = 0
+ kt2 = 3.592665704104322E-3 lkt2 = -2.007744886840338E-8 wkt2 = -1.31326041878909E-8
+ pkt2 = 7.511243690981783E-15 ua1 = 2.491910863012616E-9 lua1 = -5.539753023433691E-16
+ wua1 = 1.201122350404056E-17 pua1 = 5.425912479695583E-23 ub1 = -2.040120096307822E-18
+ lub1 = 4.127811753019636E-25 wub1 = -9.302586890018485E-26 pub1 = -9.53377561707137E-33
+ uc1 = -1.704295576853322E-10 luc1 = 6.321542381920688E-17 wuc1 = 7.969023638449497E-17
+ puc1 = -2.6240625326052E-23 at = 6.81648544644407E4 lat = 6.120169679567028E-3
+ wat = 7.282435356110214E-3 pat = -3.298095159638522E-9 prt = 0
+ njs = 1.2928 xtis = 2 tpb = 1.2287E-3
+ tpbsw = 0 tpbswg = 0 tcj = 7.92E-4
+ tcjsw = 1E-5 tcjswg = 0 tvoff = 0
+ tvfbsdoff = 0 saref = 2.74E-6 sbref = 2.74E-6
+ wlod = 0 ku0 = -2.7E-8 kvsat = 0.2
+ kvth0 = 7.9E-9 tku0 = 0 llodku0 = 0
+ wlodku0 = 1 llodvth = 0 wlodvth = 1
+ lku0 = 0 wku0 = 0 pku0 = 0
+ lkvth0 = 0 wkvth0 = 3E-7 pkvth0 = 0
+ stk2 = 0 lodk2 = 1 steta0 = 0
+ lodeta0 = 1

.model nlowvt_model.38 nmos
+ level = 54 lmin = 2.5E-7 lmax = 5E-7 wmin = 4.2E-7
+ wmax = 1E-6 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 4.148E-9
+ toxm = 4.148E-9 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 9.999999999999999E22 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {2.6E-8+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {1.2025E-8-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = -1.33E-8 dwb = -1.08E-8 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = 0.529537107912562 lvth0 = -3.563226704598899E-8
+ wvth0 = -3.217628260118897E-8 pvth0 = 4.17008003472065E-15 vfb = 0
+ k1 = 0.305576714894533 lk1 = 6.481564469523192E-8 wk1 = 4.926787199198254E-8
+ pk1 = -9.402420218106273E-15 k2 = 1.214085376494957E-3 lk2 = -1.719498935435029E-8
+ wk2 = -1.234142018909642E-8 pk2 = 2.473499960215566E-15 k3 = 1.65
+ k3b = 1.6 w0 = 1E-7 lpe0 = 2.3802E-7
+ lpeb = -4.9152E-8 vbm = -3 dvtp0 = 0
+ dvtp1 = 0 dvt0 = 0.07665 dvt1 = 0.1252
+ dvt2 = -0.05637 dvt0w = 0 dvt1w = 5.3E6
+ dvt2w = -0.032 vfbsdoff = 0 u0 = 0.023397527957844
+ lu0 = -2.295854944047906E-9 wu0 = 3.222275889747675E-9 pu0 = 2.690455976019205E-16
+ ua = -1.838712834845154E-9 lua = -1.668289468081134E-16 wua = 2.83169366621846E-16
+ pua = 1.985885945101833E-23 ub = 2.65770429695778E-18 lub = 2.15674241840549E-26
+ wub = -3.554569129997515E-26 pub = -5.190303350189236E-33 uc = 9.660112925702308E-11
+ luc = -8.305574186579605E-18 wuc = -2.497559575312107E-17 puc = 1.784464617311674E-24
+ ud = 0 up = 0 lp = 1
+ eu = 1.67 vsat = 2.640398072763062E5 lvsat = -0.024050245818725
+ wvsat = -0.068289854365778 pvsat = 1.358819414780978E-8 a0 = -0.371823946487469
+ la0 = 5.609576993606518E-7 wa0 = 8.200038294781207E-7 pa0 = -3.129732030124956E-13
+ ags = -0.490645763052312 lags = -8.160104313185405E-8 wags = 8.739018789495922E-7
+ pags = -1.500372382639959E-14 b0 = -6.087193041715727E-8 lb0 = 9.492977548555676E-15
+ wb0 = 5.77065900354651E-14 pb0 = -8.999342716030779E-21 b1 = -1.678020029772919E-9
+ lb1 = 2.616872236430865E-16 wb1 = 1.590762988224728E-15 pb1 = -2.48079488013646E-22
+ keta = 0.138212387820149 lketa = -3.436792324120019E-8 wketa = -1.078005099373271E-7
+ pketa = 2.152693162544457E-14 a1 = 0 a2 = 0.38689047
+ rdsw = 103.65 rdswmin = 0 rdw = 0
+ rdwmin = 0 rsw = 0 rswmin = 0
+ prwb = 0 prwg = 0 wr = 1
+ voff = -0.133779127377888 lvoff = 6.949674412481078E-9 wvoff = 7.816005366140176E-10
+ pvoff = -2.019350939135914E-15 voffl = 0 minv = 0
+ nfactor = 2.671625332110604 lnfactor = 2.201481799778014E-8 wnfactor = -5.532321437346928E-7
+ pnfactor = 8.427547469438754E-14 eta0 = 0.012916834918442 leta0 = -8.440057440129463E-9
+ weta0 = -9.812025035824728E-9 peta0 = 8.06594960599713E-15 etab = 8.536498091147177E-3
+ letab = -2.26559013521741E-9 wetab = -9.436980352757626E-10 petab = -1.311140607548857E-15
+ dsub = 2.437683255163648 ldsub = -4.643037106275686E-7 wdsub = -8.054533496858417E-7
+ pdsub = 1.748318921181206E-13 cit = -5.558641379310343E-6 lcit = 3.515475019655172E-12
+ wcit = 5.725580027586206E-12 pcit = -1.293694807233103E-18 cdsc = 3.8556E-37
+ cdscb = -1.1484E-4 cdscd = 4.7984E-6 pclm = 0.0384721137127
+ lpclm = 1.565953094255389E-7 wpclm = 7.105445076836033E-8 ppclm = -5.305684505905053E-14
+ pdiblc1 = 0.347645606391927 lpdiblc1 = 4.133577044179969E-8 wpdiblc1 = 4.015196514045359E-8
+ ppdiblc1 = -3.91863103788261E-14 pdiblc2 = -2.518268842261254E-3 lpdiblc2 = 3.392917318121804E-9
+ wpdiblc2 = 5.09315381590367E-9 ppdiblc2 = -1.189988636309239E-15 pdiblcb = 0
+ drout = 3.4946 pscbe1 = 4.5E8 pscbe2 = 1E-8
+ pvag = 0 delta = 0.01 fprout = 0
+ pdits = 1.4427E-15 pditsl = 0 pditsd = 0
+ lambda = 0 vtl = 0 lc = 0
+ xn = 0 alpha0 = -1.65892084510076E-3 lalpha0 = 8.473246065399912E-10
+ walpha0 = 6.138970616837762E-10 palpha0 = -2.833956995754511E-16 alpha1 = 0
+ beta0 = 18.261800506631015 lbeta0 = 3.182269325754492E-6 wbeta0 = 8.706346088153936E-7
+ pbeta0 = -7.137517610897649E-13 aigbacc = 1 bigbacc = 0
+ cigbacc = 0 nigbacc = 1 aigbinv = 0.35
+ bigbinv = 0.03 cigbinv = 6E-3 eigbinv = 1.1
+ nigbinv = 3 aigc = 0.43 bigc = 0.054
+ cigc = 0.075 aigsd = 0.43 bigsd = 0.054
+ cigsd = 0.075 dlcig = 0 nigc = 1
+ poxedge = 1 pigcd = 1 ntox = 1
+ toxref = 4.148E-9 agidl = 0 bgidl = 2.3E9
+ cgidl = 0.5 egidl = 0.8 noia = 9E41
+ noib = 1E27 noic = 8E11 em = 4.1E7
+ af = 1 ef = 1.2 kf = 0
+ lintnoi = -3E-7 tnoia = 2.5E7 tnoib = 9.9E6
+ ntnoi = 1 rnoia = 0.912 rnoib = 0.26
+ xpart = 0 cgso = {2.392894381E-10/sw_func_tox_lv_ratio} cgdo = {2.392894381E-10/sw_func_tox_lv_ratio}
+ cgbo = {1E-14/sw_func_tox_lv_ratio} ckappas = 0.6 cf = 1E-14
+ clc = 1E-7 cle = 0.6 dlc = 1.21071E-8
+ dwc = 2.6E-8 vfbcv = -1 noff = 3.8661
+ voffcv = -0.16994 acde = 0.38008 moin = 23.81
+ cgsl = {2.310725E-11/sw_func_tox_lv_ratio} cgdl = {2.310725E-11/sw_func_tox_lv_ratio} ijthsrev = 0.1
+ ijthsfwd = 0.1 xjbvs = 1 bvs = 11.9
+ jss = 2.75E-3 jsws = 6E-10 cjs = {1.210E-03*sw_func_nsd_pw_cj}
+ mjs = 0.42197 mjsws = 1E-3 cjsws = {3.230311424E-11*sw_func_nsd_pw_cj}
+ cjswgs = {1.795291232E-10*sw_func_nsd_pw_cj} mjswgs = 0.8 pbs = 0.7477
+ pbsws = 0.1 pbswgs = 0.79644 xrcrg1 = 12
+ xrcrg2 = 1 rbpb = 50 rbpd = 50
+ rbps = 50 rbdb = 50 rbsb = 50
+ gbmin = 1E-12 tnom = 30 ute = -1.419251465914213
+ lute = 1.574125181589766E-7 wute = 1.814916478466741E-7 pute = -1.047366215559618E-13
+ kt1 = -0.281105012425568 lkt1 = 1.20549038707771E-9 wkt1 = 1.035415309943829E-8
+ pkt1 = -1.36709219320369E-15 kt1l = 0 kt2 = -0.054855766789
+ lkt2 = 7.741082576689424E-9 wkt2 = 8.376418969571595E-9 pkt2 = -2.725975880812493E-15
+ ua1 = 1.262739505840201E-9 lua1 = 3.104880510284147E-17 wua1 = 4.643462829434889E-16
+ pua1 = -1.610297467432496E-22 ub1 = -1.296707708252649E-18 lub1 = 5.895404920710402E-26
+ wub1 = -3.666016277044884E-25 pub1 = 1.206746067858369E-31 uc1 = -7.636221977953907E-11
+ luc1 = 1.844407434294463E-17 wuc1 = 4.507345603516302E-17 puc1 = -9.764768718787464E-24
+ at = 1.189760600265097E5 lat = -0.0180634236077 wat = -0.011416088290731
+ pat = 5.601467170075637E-9 prt = 0 njs = 1.2928
+ xtis = 2 tpb = 1.2287E-3 tpbsw = 0
+ tpbswg = 0 tcj = 7.92E-4 tcjsw = 1E-5
+ tcjswg = 0 tvoff = 0 tvfbsdoff = 0
+ saref = 2.74E-6 sbref = 2.74E-6 wlod = 0
+ ku0 = -2.7E-8 kvsat = 0.2 kvth0 = 7.9E-9
+ tku0 = 0 llodku0 = 0 wlodku0 = 1
+ llodvth = 0 wlodvth = 1 lku0 = 0
+ wku0 = 0 pku0 = 0 lkvth0 = 0
+ wkvth0 = 3E-7 pkvth0 = 0 stk2 = 0
+ lodk2 = 1 steta0 = 0 lodeta0 = 1

.model nlowvt_model.39 nmos
+ level = 54 lmin = 1.8E-7 lmax = 2.5E-7 wmin = 4.2E-7
+ wmax = 1E-6 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 4.148E-9
+ toxm = 4.148E-9 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 9.999999999999999E22 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {2.6E-8+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {1.2025E-8-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = -1.33E-8 dwb = -1.08E-8 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = 0.736383864851615 lvth0 = -8.236929177636796E-8
+ wvth0 = -1.082958891547595E-7 pvth0 = 2.136930513549992E-14 vfb = 0
+ k1 = 0.230042524750689 lk1 = 8.188259495823346E-8 wk1 = 7.706445396491793E-8
+ pk1 = -1.568305791489102E-14 k2 = 0.02437038930911 lk2 = -2.242715622792469E-8
+ wk2 = -2.086294003629927E-8 pk2 = 4.398937369691051E-15 k3 = 1.65
+ k3b = 1.6 w0 = 1E-7 lpe0 = 2.3802E-7
+ lpeb = -4.9152E-8 vbm = -3 dvtp0 = 0
+ dvtp1 = 0 dvt0 = 0.07665 dvt1 = 0.1252
+ dvt2 = -0.05637 dvt0w = 0 dvt1w = 5.3E6
+ dvt2w = -0.032 vfbsdoff = 0 u0 = 0.021731413379893
+ lu0 = -1.919396355159838E-9 wu0 = 3.83540605443282E-9 pu0 = 1.30508836891312E-16
+ ua = -2.612753463107833E-9 lua = 8.06553314783895E-18 wua = 5.680163178225121E-16
+ pua = -4.450230917277218E-23 ub = 3.607558224297483E-18 lub = -1.930520706983512E-25
+ wub = -3.850919365609857E-25 pub = 7.378967076653609E-32 uc = 9.008944408093003E-11
+ luc = -6.834258921041383E-18 wuc = -2.257929560831883E-17 puc = 1.243020599593608E-24
+ ud = 0 up = 0 lp = 1
+ eu = 1.67 vsat = 1.525062300050906E5 lvsat = 1.150765965706118E-3
+ wvsat = -0.027245497929969 pvsat = 4.314221811138631E-9 a0 = 6.813486837882976
+ la0 = -1.06256327236785E-6 wa0 = -1.824190539170204E-6 pa0 = 2.844825145835932E-13
+ ags = -5.180926930301574 lags = 9.781679866081169E-7 wags = 2.599925348497321E-6
+ pags = -4.04998726770709E-13 b0 = -6.087193041715728E-8 lb0 = 9.492977548555682E-15
+ wb0 = 5.770659003546511E-14 pb0 = -8.999342716030784E-21 b1 = -1.678020029772924E-9
+ lb1 = 2.616872236430874E-16 wb1 = 1.590762988224731E-15 pb1 = -2.480794880136468E-22
+ keta = 0.329834310725622 lketa = -7.766489672169184E-8 wketa = -1.783173775665414E-7
+ pketa = 3.746021786626555E-14 a1 = 0 a2 = 0.38689047
+ rdsw = 103.65 rdswmin = 0 rdw = 0
+ rdwmin = 0 rsw = 0 rswmin = 0
+ prwb = 0 prwg = 0 wr = 1
+ voff = -0.184998766545315 lvoff = 1.852275188236126E-8 wvoff = 1.963042775022762E-8
+ pvoff = -6.278243448051905E-15 voffl = 0 minv = 0
+ nfactor = 1.167837466878308 lnfactor = 3.617956861470175E-7 wnfactor = 1.617906707926484E-10
+ pnfactor = -4.076388478453188E-14 eta0 = -0.24694514621595 leta0 = 5.02757571971863E-8
+ weta0 = 8.581718402163191E-8 peta0 = -1.354147018053519E-14 etab = 0.023576290085277
+ letab = -5.663831136290958E-9 wetab = -6.478341489115669E-9 petab = -6.058791915373025E-17
+ dsub = 0.451152321508408 ldsub = -1.54470461681673E-8 wdsub = -7.440996610071383E-8
+ pdsub = 9.652639597060944E-15 cit = 2.820697044334976E-5 lcit = -4.113864971674879E-12
+ wcit = -6.700165123152715E-12 pcit = 1.513902309576356E-18 cdsc = 3.8556E-37
+ cdscb = -1.1484E-4 cdscd = 4.7984E-6 pclm = 1.914566679383637
+ lpclm = -2.673082576878092E-7 wpclm = -6.193483493985449E-7 ppclm = 1.029396676386617E-13
+ pdiblc1 = -1.873604787696745 lpdiblc1 = 5.432272969861349E-7 wpdiblc1 = 8.575721101650849E-7
+ ppdiblc1 = -2.238823921471415E-13 pdiblc2 = 5.341922794666685E-3 lpdiblc2 = 1.616907017757937E-9
+ wpdiblc2 = 2.200603293513125E-9 ppdiblc2 = -5.364168457750959E-16 pdiblcb = 0
+ drout = 3.4946 pscbe1 = 4.5E8 pscbe2 = 1E-8
+ pvag = 0 delta = 0.01 fprout = 0
+ pdits = 1.4427E-15 pditsl = 0 pditsd = 0
+ lambda = 0 vtl = 0 lc = 0
+ xn = 0 alpha0 = 5.743735433277913E-3 lalpha0 = -8.253055795596699E-10
+ walpha0 = -2.110280448759576E-9 palpha0 = 3.321322089092242E-16 alpha1 = 0
+ beta0 = 41.622826806308055 lbeta0 = -2.096154566657535E-6 wbeta0 = -7.726223069465755E-6
+ pbeta0 = 1.22870823131786E-12 aigbacc = 1 bigbacc = 0
+ cigbacc = 0 nigbacc = 1 aigbinv = 0.35
+ bigbinv = 0.03 cigbinv = 6E-3 eigbinv = 1.1
+ nigbinv = 3 aigc = 0.43 bigc = 0.054
+ cigc = 0.075 aigsd = 0.43 bigsd = 0.054
+ cigsd = 0.075 dlcig = 0 nigc = 1
+ poxedge = 1 pigcd = 1 ntox = 1
+ toxref = 4.148E-9 agidl = 0 bgidl = 2.3E9
+ cgidl = 0.5 egidl = 0.8 noia = 9E41
+ noib = 1E27 noic = 8E11 em = 4.1E7
+ af = 1 ef = 1.2 kf = 0
+ lintnoi = -3E-7 tnoia = 2.5E7 tnoib = 9.9E6
+ ntnoi = 1 rnoia = 0.912 rnoib = 0.26
+ xpart = 0 cgso = {2.392894381E-10/sw_func_tox_lv_ratio} cgdo = {2.392894381E-10/sw_func_tox_lv_ratio}
+ cgbo = {1E-14/sw_func_tox_lv_ratio} ckappas = 0.6 cf = 1E-14
+ clc = 1E-7 cle = 0.6 dlc = 1.21071E-8
+ dwc = 2.6E-8 vfbcv = -1 noff = 3.8661
+ voffcv = -0.16994 acde = 0.38008 moin = 23.81
+ cgsl = {2.310725E-11/sw_func_tox_lv_ratio} cgdl = {2.310725E-11/sw_func_tox_lv_ratio} ijthsrev = 0.1
+ ijthsfwd = 0.1 xjbvs = 1 bvs = 11.9
+ jss = 2.75E-3 jsws = 6E-10 cjs = {1.210E-03*sw_func_nsd_pw_cj}
+ mjs = 0.42197 mjsws = 1E-3 cjsws = {3.230311424E-11*sw_func_nsd_pw_cj}
+ cjswgs = {1.795291232E-10*sw_func_nsd_pw_cj} mjswgs = 0.8 pbs = 0.7477
+ pbsws = 0.1 pbswgs = 0.79644 xrcrg1 = 12
+ xrcrg2 = 1 rbpb = 50 rbpd = 50
+ rbps = 50 rbdb = 50 rbsb = 50
+ gbmin = 1E-12 tnom = 30 ute = 1.612684878144899
+ lute = -5.276534987811798E-7 wute = -9.34260926767078E-7 pute = 1.473676726780155E-13
+ kt1 = -0.162832527755616 lkt1 = -2.55181775240979E-8 wkt1 = -3.317012125910475E-8
+ pkt1 = 8.467217598109107E-15 kt1l = 0 kt2 = -0.032869986014417
+ lkt2 = 2.773395410672422E-9 wkt2 = 2.856516445241667E-10 pkt2 = -8.978670037180266E-16
+ ua1 = 5.271837688854984E-9 lua1 = -8.748069293493484E-16 wua1 = -1.011001848405952E-15
+ pua1 = 1.723251635351564E-22 ub1 = -4.690881959509792E-18 lub1 = 8.258677212786556E-25
+ wub1 = 8.824544967581407E-25 pub1 = -1.615496245364941E-31 uc1 = -3.005290485666221E-11
+ luc1 = 7.980484636120608E-18 wuc1 = 2.803162814354433E-17 puc1 = -5.91416770667622E-24
+ at = -4.503950501309626E4 lat = 0.018995893312999 wat = 0.048941639643844
+ pat = -8.036361456741578E-9 prt = 0 njs = 1.2928
+ xtis = 2 tpb = 1.2287E-3 tpbsw = 0
+ tpbswg = 0 tcj = 7.92E-4 tcjsw = 1E-5
+ tcjswg = 0 tvoff = 0 tvfbsdoff = 0
+ saref = 2.74E-6 sbref = 2.74E-6 wlod = 0
+ ku0 = -2.7E-8 kvsat = 0.2 kvth0 = 7.9E-9
+ tku0 = 0 llodku0 = 0 wlodku0 = 1
+ llodvth = 0 wlodvth = 1 lku0 = 0
+ wku0 = 0 pku0 = 0 lkvth0 = 0
+ wkvth0 = 3E-7 pkvth0 = 0 stk2 = 0
+ lodk2 = 1 steta0 = 0 lodeta0 = 1

.model nlowvt_model.40 nmos
+ level = 54 lmin = 1.5E-7 lmax = 1.8E-7 wmin = 4.2E-7
+ wmax = 1E-6 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 4.148E-9
+ toxm = 4.148E-9 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 9.999999999999999E22 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {2.6E-8+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {1.2025E-8-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = -1.33E-8 dwb = -1.08E-8 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = -0.260340008328966 lvth0 = 7.306979624614356E-8
+ wvth0 = 3.482045360250594E-7 pvth0 = -4.982193617129284E-14 vfb = 0
+ k1 = 1.291281131149425 lk1 = -8.361756570964946E-8 wk1 = -2.623134781296553E-7
+ pk1 = 3.724293059525767E-14 k2 = -0.259338002614104 lk2 = 2.181716749250047E-8
+ wk2 = 4.665847916759008E-8 pk2 = -6.131027955155493E-15 k3 = 1.65
+ k3b = 1.6 w0 = 1E-7 lpe0 = 2.3802E-7
+ lpeb = -4.9152E-8 vbm = -3 dvtp0 = 0
+ dvtp1 = 0 dvt0 = 0.07665 dvt1 = 0.1252
+ dvt2 = -0.05637 dvt0w = 0 dvt1w = 5.3E6
+ dvt2w = -0.032 vfbsdoff = 0 u0 = -0.031789832207931
+ lu0 = 6.427241894261327E-9 wu0 = 3.297514022531862E-8 pu0 = -4.413832707058328E-15
+ ua = -4.860133603401842E-9 lua = 3.585444660266894E-16 wua = 1.848748842574544E-15
+ pua = -2.442325464078515E-22 ub = 2.51336711674069E-18 lub = -2.241296747486911E-26
+ wub = 1.451323821594265E-25 pub = -8.898811737912189E-33 uc = 1.871521082712311E-10
+ luc = -2.197118140151883E-17 wuc = -6.382021977981304E-17 puc = 7.674542724138128E-24
+ ud = 0 up = 0 lp = 1
+ eu = 1.67 vsat = 1.588356211183908E5 lvsat = 1.63697421586955E-4
+ wvsat = 8.187328417765502E-3 pvsat = -1.21152745779053E-9 a0 = 0
+ ags = 0.435938548275863 lags = 1.022178152239654E-7 wags = 2.213923023448227E-8
+ pags = -2.992981627619243E-15 b0 = 0 b1 = 0
+ keta = -1.224127403398735 lketa = 1.646754325960018E-7 wketa = 6.534128831174013E-7
+ pketa = -9.224811628739532E-14 a1 = 0 a2 = 0.38689047
+ rdsw = 103.65 rdswmin = 0 rdw = 0
+ rdwmin = 0 rsw = 0 rswmin = 0
+ prwb = 0 prwg = 0 wr = 1
+ voff = 0.210568999513494 lvoff = -4.316604123451014E-8 wvoff = -1.837892608759526E-7
+ pvoff = 2.54450569932009E-14 voffl = 0 minv = 0
+ nfactor = 4.594499715021837 lnfactor = -1.725922914509658E-7 wnfactor = -1.862683961546702E-6
+ pnfactor = 2.497469102737864E-13 eta0 = 0.140369114003425 leta0 = -1.012590168402521E-8
+ weta0 = 4.230789679767283E-8 peta0 = -6.756196837958777E-15 etab = 8.421899546183914E-3
+ letab = -3.300503931719449E-9 wetab = -5.996617802294236E-8 petab = 8.28084018829654E-15
+ dsub = 0.738875246707356 ldsub = -6.031743635294325E-8 wdsub = -6.515108323097376E-8
+ pdsub = 8.208716813524979E-15 cit = -3.248293103448277E-5 lcit = 5.350725163793104E-12
+ wcit = 1.563371862068966E-11 pcit = -1.969066860275862E-18 cdsc = 3.8556E-37
+ cdscb = -1.1484E-4 cdscd = 4.7984E-6 pclm = -0.249078158505747
+ lpclm = 7.011215478104019E-8 wpclm = 1.211117164634482E-7 ppclm = -1.253507963251613E-14
+ pdiblc1 = 4.512860269409426 lpdiblc1 = -4.527419286695723E-7 wpdiblc1 = -3.131112765809336E-6
+ ppdiblc1 = 3.981530142610693E-13 pdiblc2 = 0.061154042401149 lpdiblc2 = -7.086993034873044E-9
+ wpdiblc2 = -1.699993691028965E-8 ppdiblc2 = 2.457907399007947E-15 pdiblcb = 0
+ drout = 3.4946 pscbe1 = 4.5E8 pscbe2 = 1E-8
+ pvag = 0 delta = 0.01 fprout = 0
+ pdits = 1.4427E-15 pditsl = 0 pditsd = 0
+ lambda = 0 vtl = 0 lc = 0
+ xn = 0 alpha0 = 1.410962310681609E-3 lalpha0 = -1.496096110907762E-10
+ walpha0 = 2.496919155942347E-10 palpha0 = -3.590548131175251E-17 alpha1 = 0
+ beta0 = 32.16213007719541 lbeta0 = -6.207589117524169E-7 wbeta0 = 2.176484219138757E-6
+ pbeta0 = -3.156189703400131E-13 aigbacc = 1 bigbacc = 0
+ cigbacc = 0 nigbacc = 1 aigbinv = 0.35
+ bigbinv = 0.03 cigbinv = 6E-3 eigbinv = 1.1
+ nigbinv = 3 aigc = 0.43 bigc = 0.054
+ cigc = 0.075 aigsd = 0.43 bigsd = 0.054
+ cigsd = 0.075 dlcig = 0 nigc = 1
+ poxedge = 1 pigcd = 1 ntox = 1
+ toxref = 4.148E-9 agidl = 0 bgidl = 2.3E9
+ cgidl = 0.5 egidl = 0.8 noia = 9E41
+ noib = 1E27 noic = 8E11 em = 4.1E7
+ af = 1 ef = 1.2 kf = 0
+ lintnoi = -3E-7 tnoia = 2.5E7 tnoib = 9.9E6
+ ntnoi = 1 rnoia = 0.912 rnoib = 0.26
+ xpart = 0 cgso = {2.392894381E-10/sw_func_tox_lv_ratio} cgdo = {2.392894381E-10/sw_func_tox_lv_ratio}
+ cgbo = {1E-14/sw_func_tox_lv_ratio} ckappas = 0.6 cf = 1E-14
+ clc = 1E-7 cle = 0.6 dlc = 1.21071E-8
+ dwc = 2.6E-8 vfbcv = -1 noff = 3.8661
+ voffcv = -0.16994 acde = 0.38008 moin = 23.81
+ cgsl = {2.310725E-11/sw_func_tox_lv_ratio} cgdl = {2.310725E-11/sw_func_tox_lv_ratio} ijthsrev = 0.1
+ ijthsfwd = 0.1 xjbvs = 1 bvs = 11.9
+ jss = 2.75E-3 jsws = 6E-10 cjs = {1.210E-03*sw_func_nsd_pw_cj}
+ mjs = 0.42197 mjsws = 1E-3 cjsws = {3.230311424E-11*sw_func_nsd_pw_cj}
+ cjswgs = {1.795291232E-10*sw_func_nsd_pw_cj} mjswgs = 0.8 pbs = 0.7477
+ pbsws = 0.1 pbswgs = 0.79644 xrcrg1 = 12
+ xrcrg2 = 1 rbpb = 50 rbpd = 50
+ rbps = 50 rbdb = 50 rbsb = 50
+ gbmin = 1E-12 tnom = 30 ute = -2.445538344827586
+ lute = 1.052264128413792E-7 wute = 2.316662468965515E-7 pute = -3.445867005482755E-14
+ kt1 = -0.531037394367816 lkt1 = 3.190337142407469E-8 wkt1 = 1.709223880606896E-7
+ pkt1 = -2.336100923031282E-14 kt1l = 0 kt2 = -0.075960689968966
+ lkt2 = 9.493390692384315E-9 wkt2 = 7.633534285793268E-10 pkt2 = -9.723645969414283E-16
+ ua1 = -1.599231564712644E-9 lua1 = 1.96736320744523E-16 wua1 = 7.822840523475864E-16
+ pua1 = -1.073377726873578E-22 ub1 = 1.49963842137931E-18 lub1 = -1.395439321209999E-25
+ wub1 = -7.305231006675861E-25 pub1 = 8.999423178204797E-32 uc1 = 2.503911781931034E-10
+ luc1 = -3.575477011549034E-17 wuc1 = -1.325399130470621E-16 puc1 = 1.912696414199884E-23
+ at = 9.111705956321838E4 lat = -2.237722932677011E-3 wat = -0.015213759545931
+ pat = 1.968673046903807E-9 prt = 0 njs = 1.2928
+ xtis = 2 tpb = 1.2287E-3 tpbsw = 0
+ tpbswg = 0 tcj = 7.92E-4 tcjsw = 1E-5
+ tcjswg = 0 tvoff = 0 tvfbsdoff = 0
+ saref = 1.1E-6 sbref = 1.1E-6 wlod = 0
+ ku0 = -2.7E-8 kvsat = 0.2 kvth0 = 7.9E-9
+ tku0 = 0 llodku0 = 0 wlodku0 = 1
+ llodvth = 0 wlodvth = 1 lku0 = 0
+ wku0 = 0 pku0 = 0 lkvth0 = 0
+ wkvth0 = 3E-7 pkvth0 = 0 stk2 = 0
+ lodk2 = 1 steta0 = 0 lodeta0 = 1

.ends sky130_fd_pr__nfet_01v8_lvt
