* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

******************************************************************
******************************************************************
*  *****************************************************
*  12/08/2020 Usman Suriono
*      Why     : New scalable sky130_fd_pr__nfet_01v8 5V (HV) model
*      What    : Converted from discrete nhv models
*                Replaced rsh from 1 to calculated rsh from the original model.
*                PDK netlist nrd/nrs = ratio of distance the middle of the contact to Gate.
*
*  *****************************************************
*
*  Nmos HV 5V Model
*  -----------------------------------------------------

.subckt  sky130_fd_pr__nfet_g5v0d10v5  d g s b  mult=1
+ 
.param  l = 1 w = 1 nf = 1 ad = 0 as = 0 pd = 0 ps = 0 nrd = {0.14/w} nrs = {0.14/w} sa = 0 sb = 0 sd = 0
+ swx_nrds = {89.1*nf/w+443.5}
+ swx_vth = {sw_vth0_sky130_fd_pr__nfet_g5v0d10v5+sw_vth0_sky130_fd_pr__nfet_g5v0d10v5_mc}

Msky130_fd_pr__nfet_g5v0d10v5  d g s b nhv_model l = {l} w = {w} ad = {ad} as = {as} pd = {pd} ps = {ps} nrd = {nrd} nrs = {nrs} sa = {sa} sb = {sb} sd = {sd} nf = {nf}
* + deltox = 0.3*(sw_tox_hv_corner - sw_tox_hv_nom) + sw_tox_hv_mc + sw_mm_tox_hv * mismatch_factor*MC_MM_SWITCH*AGAUSS(0,1.0,1)/sqrt(l*w*mult)
* + mulu0  = sw_u0_sky130_fd_pr__nfet_g5v0d10v5
+ delvto = {swx_vth*(0.10*8/l+0.90)*(0.045*7/w+0.955)*(-0.0007*56/(l*w)+1.0007)+sw_mm_vth0_sky130_fd_pr__nfet_g5v0d10v5*mismatch_factor*MC_MM_SWITCH*AGAUSS(0,1.0,1)/sqrt(l*w*mult)}
* + mulvsat = sw_vsat_sky130_fd_pr__nfet_g5v0d10v5




.model nhv_model.1 nmos
+ level = 54 lmin = 8E-6 lmax = 2.02E-5 wmin = 2E-5
+ wmax = 1.01E-3 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 1.16E-8
+ toxm = 1.16E-8 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 1E23 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {2.1346E-8+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {7.6507E-8-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = -4.1292E-9 dwb = -1.6944E-9 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = 0.78882 k1 = 0.88325
+ k2 = -0.039667 k3 = -0.884 k3b = 0.43
+ w0 = 0 lpe0 = 2.5E-8 lpeb = -2.182E-7
+ vbm = -3 dvtp0 = 0 dvtp1 = 0
+ dvt0 = 0 dvt1 = 0.53 dvt2 = -0.19251
+ dvt0w = 0.16 dvt1w = 6.9091E6 dvt2w = -0.036016
+ vfbsdoff = 0 u0 = 4.21082E-2 ua = -5.92431E-11
+ ub = 1.71671E-18 uc = 6.6204E-11 ud = 0
+ up = 0 lp = 1 eu = 1.67
+ vsat = 1.0566E5 a0 = 0.942599 ags = 0.149418
+ b0 = 3.2933E-8 b1 = 0 keta = -0.02132
+ a1 = 0 a2 = 0.659726 rdsw = 724.62
+ rdswmin = 0 rdw = 0 rdwmin = 0
+ rsw = 0 rswmin = 0 prwb = 0.05626
+ prwg = 0.048 wr = 1 voff = -0.20613
+ voffl = -4.257949E-7 minv = 0 nfactor = 0.96538
+ eta0 = 0.032 etab = -0.01932 dsub = 0.504
+ cit = -8E-4 cdsc = 0 cdscb = 0
+ cdscd = 0 pclm = 0.33405 pdiblc1 = 0.21098
+ pdiblc2 = 2E-4 pdiblcb = -0.26831 drout = 0.36075
+ pscbe1 = 9.3731E8 pscbe2 = 1.68E-6 pvag = 1.99
+ delta = 0.0246 fprout = 10.125 pdits = 0
+ pditsl = 0 pditsd = 0 lambda = 0
+ vtl = 0 lc = 5E-9 xn = 3
+ alpha0 = 1.4467E-5 alpha1 = 0 beta0 = 24
+ aigbacc = 1 bigbacc = 0 cigbacc = 0
+ nigbacc = 1 aigbinv = 0.35 bigbinv = 0.03
+ cigbinv = 6E-3 eigbinv = 1.1 nigbinv = 3
+ aigc = 0.43 bigc = 0.054 cigc = 0.075
+ aigsd = 0.43 bigsd = 0.054 cigsd = 0.075
+ dlcig = 0 nigc = 1 poxedge = 1
+ pigcd = 1 ntox = 1 toxref = 1.16E-8
+ agidl = 5.06E-11 bgidl = 1.058E9 cgidl = 4E3
+ egidl = 0.8 noia = 2.6E41 noib = 0
+ noic = 0 em = 4.1E7 af = 1
+ ef = 0.89 kf = 0 lintnoi = 0
+ tnoia = 7.5E6 tnoib = 7.2E6 ntnoi = 1
+ rnoia = 0.794 rnoib = 0.38 xpart = 0
+ cgso = {2.754679E-10/sw_func_tox_hv_ratio} cgdo = {2.754679E-10/sw_func_tox_hv_ratio} cgbo = {0/sw_func_tox_hv_ratio}
+ ckappas = 0.6 cf = 0 clc = 1E-7
+ cle = 0.6 dlc = 6.5995E-8 dwc = 0
+ vfbcv = -1 noff = 4 voffcv = -0.4104
+ acde = 0.4176 moin = 15 cgsl = {4.49025E-11/sw_func_tox_hv_ratio}
+ cgdl = {4.49025E-11/sw_func_tox_hv_ratio} ijthsrev = 0.1 ijthsfwd = 0.1
+ xjbvs = 1 bvs = 12.636 jss = 3.75E-4
+ jsws = 5.84E-11 cjs = {8.310E-04*sw_func_nsd_pw_cj} mjs = 0.295
+ mjsws = 0.037586 cjsws = {8.643094E-11*sw_func_nsd_pw_cj} cjswgs = {5.47776E-11*sw_func_nsd_pw_cj}
+ mjswgs = 0.78692 pbs = 0.72468 pbsws = 0.29067
+ pbswgs = 0.54958 xrcrg1 = 12 xrcrg2 = 1
+ rbpb = 50 rbpd = 50 rbps = 50
+ rbdb = 50 rbsb = 50 gbmin = 1E-12
+ tnom = 30 ute = -1.2986 kt1 = -0.40273
+ kt1l = 0 kt2 = -0.019151 ua1 = 3.0044E-9
+ ub1 = -3.7525E-18 uc1 = -5.9821E-11 at = 1.6E5
+ prt = 0 njs = 1.0773 xtis = 0.76
+ tpb = 1.344E-3 tpbsw = 9.9005E-4 tpbswg = 0
+ tcj = 6.7434E-4 tcjsw = 2.493E-4 tcjswg = 0
+ tvoff = 0 tvfbsdoff = 0 saref = 3E-6
+ sbref = 3E-6 wlod = 0 ku0 = -4.5E-8
+ kvsat = 0.3 kvth0 = 1.1E-8 tku0 = 0
+ llodku0 = 0 wlodku0 = 1 llodvth = 0
+ wlodvth = 1 lku0 = 0 wku0 = 2E-7
+ pku0 = 0 lkvth0 = 0 wkvth0 = 6.5E-7
+ pkvth0 = 0 stk2 = 0 lodk2 = 1
+ steta0 = 0 lodeta0 = 1

.model nhv_model.2 nmos
+ level = 54 lmin = 4E-6 lmax = 8E-6 wmin = 2E-5
+ wmax = 1.01E-3 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 1.16E-8
+ toxm = 1.16E-8 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 1E23 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {2.1346E-8+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {7.6507E-8-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = -4.1292E-9 dwb = -1.6944E-9 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = 0.783367 lvth0 = 4.279042E-8
+ k1 = 0.88325 k2 = -4.10016E-2 lk2 = 1.047271E-8
+ k3 = -0.884 k3b = 0.43 w0 = 0
+ lpe0 = 2.5E-8 lpeb = -2.182E-7 vbm = -3
+ dvtp0 = 0 dvtp1 = 0 dvt0 = 0
+ dvt1 = 0.53 dvt2 = -0.19251 dvt0w = 0.16
+ dvt1w = 6.9091E6 dvt2w = -0.036016 vfbsdoff = 0
+ u0 = 4.15573E-2 lu0 = 4.322814E-9 ua = -1.016037E-10
+ lua = 3.324031E-16 ub = 1.752362E-18 lub = -2.797603E-25
+ uc = 6.6204E-11 ud = 0 up = 0
+ lp = 1 eu = 1.67 vsat = 1.104687E5
+ lvsat = -3.77341E-2 a0 = 1.033611 la0 = -7.141721E-7
+ ags = 0.152066 lags = -2.078241E-8 b0 = 3.2933E-8
+ b1 = 0 keta = -1.72682E-2 lketa = -3.179472E-8
+ a1 = 0 a2 = 0.659726 rdsw = 724.62
+ rdswmin = 0 rdw = 0 rdwmin = 0
+ rsw = 0 rswmin = 0 prwb = 0.05626
+ prwg = 0.048 wr = 1 voff = -0.20613
+ voffl = -4.257949E-7 minv = 0 nfactor = 1.012092
+ lnfactor = -3.665486E-7 eta0 = 0.032 etab = -0.01932
+ dsub = 0.504 cit = -8E-4 cdsc = 0
+ cdscb = 0 cdscd = 0 pclm = 0.259909
+ lpclm = 5.817837E-7 pdiblc1 = 0.21098 pdiblc2 = 2E-4
+ pdiblcb = -0.26831 drout = 0.36075 pscbe1 = 9.3731E8
+ pscbe2 = 1.68E-6 pvag = 1.99 delta = 0.0246
+ fprout = 10.125 pdits = 0 pditsl = 0
+ pditsd = 0 lambda = 0 vtl = 0
+ lc = 5E-9 xn = 3 alpha0 = 1.4467E-5
+ alpha1 = 0 beta0 = 21.499459 lbeta0 = 1.962171E-5
+ aigbacc = 1 bigbacc = 0 cigbacc = 0
+ nigbacc = 1 aigbinv = 0.35 bigbinv = 0.03
+ cigbinv = 6E-3 eigbinv = 1.1 nigbinv = 3
+ aigc = 0.43 bigc = 0.054 cigc = 0.075
+ aigsd = 0.43 bigsd = 0.054 cigsd = 0.075
+ dlcig = 0 nigc = 1 poxedge = 1
+ pigcd = 1 ntox = 1 toxref = 1.16E-8
+ agidl = 5.06E-11 bgidl = 1.058E9 cgidl = 4E3
+ egidl = 0.8 noia = 2.6E41 noib = 0
+ noic = 0 em = 4.1E7 af = 1
+ ef = 0.89 kf = 0 lintnoi = 0
+ tnoia = 7.5E6 tnoib = 7.2E6 ntnoi = 1
+ rnoia = 0.794 rnoib = 0.38 xpart = 0
+ cgso = {2.754679E-10/sw_func_tox_hv_ratio} cgdo = {2.754679E-10/sw_func_tox_hv_ratio} cgbo = {0/sw_func_tox_hv_ratio}
+ ckappas = 0.6 cf = 0 clc = 1E-7
+ cle = 0.6 dlc = 6.5995E-8 dwc = 0
+ vfbcv = -1 noff = 4 voffcv = -0.4104
+ acde = 0.4176 moin = 15 cgsl = {4.49025E-11/sw_func_tox_hv_ratio}
+ cgdl = {4.49025E-11/sw_func_tox_hv_ratio} ijthsrev = 0.1 ijthsfwd = 0.1
+ xjbvs = 1 bvs = 12.636 jss = 3.75E-4
+ jsws = 5.84E-11 cjs = {8.310E-04*sw_func_nsd_pw_cj} mjs = 0.295
+ mjsws = 0.037586 cjsws = {8.643094E-11*sw_func_nsd_pw_cj} cjswgs = {5.47776E-11*sw_func_nsd_pw_cj}
+ mjswgs = 0.78692 pbs = 0.72468 pbsws = 0.29067
+ pbswgs = 0.54958 xrcrg1 = 12 xrcrg2 = 1
+ rbpb = 50 rbpd = 50 rbps = 50
+ rbdb = 50 rbsb = 50 gbmin = 1E-12
+ tnom = 30 ute = -1.33707 lute = 3.018725E-7
+ kt1 = -0.414271 lkt1 = 9.056174E-8 kt1l = 0
+ kt2 = -0.019151 ua1 = 3.0044E-9 ub1 = -3.7525E-18
+ uc1 = -5.9821E-11 at = 2.369397E5 lat = -0.603745
+ prt = 0 njs = 1.0773 xtis = 0.76
+ tpb = 1.344E-3 tpbsw = 9.9005E-4 tpbswg = 0
+ tcj = 6.7434E-4 tcjsw = 2.493E-4 tcjswg = 0
+ tvoff = 0 tvfbsdoff = 0 saref = 3E-6
+ sbref = 3E-6 wlod = 0 ku0 = -4.5E-8
+ kvsat = 0.3 kvth0 = 1.1E-8 tku0 = 0
+ llodku0 = 0 wlodku0 = 1 llodvth = 0
+ wlodvth = 1 lku0 = 0 wku0 = 2E-7
+ pku0 = 0 lkvth0 = 0 wkvth0 = 6.5E-7
+ pkvth0 = 0 stk2 = 0 lodk2 = 1
+ steta0 = 0 lodeta0 = 1

.model nhv_model.3 nmos
+ level = 54 lmin = 2E-6 lmax = 4E-6 wmin = 2E-5
+ wmax = 1.01E-3 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 1.16E-8
+ toxm = 1.16E-8 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 1E23 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {2.1346E-8+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {7.6507E-8-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = -4.1292E-9 dwb = -1.6944E-9 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = 0.799231 lvth0 = -1.823938E-8
+ k1 = 0.88325 k2 = -4.25688E-2 lk2 = 1.650177E-8
+ k3 = -0.884 k3b = 0.43 w0 = 0
+ lpe0 = 2.5E-8 lpeb = -2.182E-7 vbm = -3
+ dvtp0 = 0 dvtp1 = 0 dvt0 = 0
+ dvt1 = 0.53 dvt2 = -0.19251 dvt0w = 0.16
+ dvt1w = 6.9091E6 dvt2w = -0.036016 vfbsdoff = 0
+ u0 = 4.27638E-2 lu0 = -3.18674E-10 ua = 1.059937E-10
+ lua = -4.662212E-16 ub = 1.549686E-18 lub = 4.99931E-25
+ uc = 6.6204E-11 ud = 0 up = 0
+ lp = 1 eu = 1.67 vsat = 9.377998E4
+ lvsat = 2.64674E-2 a0 = 0.476534 la0 = 1.428898E-6
+ ags = 0.119435 lags = 1.047503E-7 b0 = 3.2933E-8
+ b1 = 0 keta = -3.92681E-2 lketa = 5.283878E-8
+ a1 = 0 a2 = 0.659726 rdsw = 724.62
+ rdswmin = 0 rdw = 0 rdwmin = 0
+ rsw = 0 rswmin = 0 prwb = 0.05626
+ prwg = 0.048 wr = 1 voff = -0.20613
+ voffl = -4.257949E-7 minv = 0 nfactor = 0.961332
+ lnfactor = -1.71274E-7 eta0 = 0.032 etab = -0.01932
+ dsub = 0.504 cit = -8E-4 cdsc = 0
+ cdscb = 0 cdscd = 0 pclm = 0.600982
+ lpclm = -7.303213E-7 pdiblc1 = 0.21098 pdiblc2 = 2E-4
+ pdiblcb = -0.26831 drout = 0.36075 pscbe1 = 9.3731E8
+ pscbe2 = 1.68E-6 pvag = 1.99 delta = 0.0246
+ fprout = 10.125 pdits = 0 pditsl = 0
+ pditsd = 0 lambda = 0 vtl = 0
+ lc = 5E-9 xn = 3 alpha0 = 1.4467E-5
+ alpha1 = 0 beta0 = 23.859073 lbeta0 = 1.054431E-5
+ aigbacc = 1 bigbacc = 0 cigbacc = 0
+ nigbacc = 1 aigbinv = 0.35 bigbinv = 0.03
+ cigbinv = 6E-3 eigbinv = 1.1 nigbinv = 3
+ aigc = 0.43 bigc = 0.054 cigc = 0.075
+ aigsd = 0.43 bigsd = 0.054 cigsd = 0.075
+ dlcig = 0 nigc = 1 poxedge = 1
+ pigcd = 1 ntox = 1 toxref = 1.16E-8
+ agidl = 5.06E-11 bgidl = 1.058E9 cgidl = 4E3
+ egidl = 0.8 noia = 2.6E41 noib = 0
+ noic = 0 em = 4.1E7 af = 1
+ ef = 0.89 kf = 0 lintnoi = 0
+ tnoia = 7.5E6 tnoib = 7.2E6 ntnoi = 1
+ rnoia = 0.794 rnoib = 0.38 xpart = 0
+ cgso = {2.754679E-10/sw_func_tox_hv_ratio} cgdo = {2.754679E-10/sw_func_tox_hv_ratio} cgbo = {0/sw_func_tox_hv_ratio}
+ ckappas = 0.6 cf = 0 clc = 1E-7
+ cle = 0.6 dlc = 6.5995E-8 dwc = 0
+ vfbcv = -1 noff = 4 voffcv = -0.4104
+ acde = 0.4176 moin = 15 cgsl = {4.49025E-11/sw_func_tox_hv_ratio}
+ cgdl = {4.49025E-11/sw_func_tox_hv_ratio} ijthsrev = 0.1 ijthsfwd = 0.1
+ xjbvs = 1 bvs = 12.636 jss = 3.75E-4
+ jsws = 5.84E-11 cjs = {8.310E-04*sw_func_nsd_pw_cj} mjs = 0.295
+ mjsws = 0.037586 cjsws = {8.643094E-11*sw_func_nsd_pw_cj} cjswgs = {5.47776E-11*sw_func_nsd_pw_cj}
+ mjswgs = 0.78692 pbs = 0.72468 pbsws = 0.29067
+ pbswgs = 0.54958 xrcrg1 = 12 xrcrg2 = 1
+ rbpb = 50 rbpd = 50 rbps = 50
+ rbdb = 50 rbsb = 50 gbmin = 1E-12
+ tnom = 30 ute = -1.22166 lute = -1.421066E-7
+ kt1 = -0.407353 lkt1 = 6.394796E-8 kt1l = 0
+ kt2 = -0.019151 ua1 = 3.0044E-9 ub1 = -3.7525E-18
+ uc1 = -5.9821E-11 at = 1.391036E5 lat = -0.227371
+ prt = 0 njs = 1.0773 xtis = 0.76
+ tpb = 1.344E-3 tpbsw = 9.9005E-4 tpbswg = 0
+ tcj = 6.7434E-4 tcjsw = 2.493E-4 tcjswg = 0
+ tvoff = 0 tvfbsdoff = 0 saref = 3E-6
+ sbref = 3E-6 wlod = 0 ku0 = -4.5E-8
+ kvsat = 0.3 kvth0 = 1.1E-8 tku0 = 0
+ llodku0 = 0 wlodku0 = 1 llodvth = 0
+ wlodvth = 1 lku0 = 0 wku0 = 2E-7
+ pku0 = 0 lkvth0 = 0 wkvth0 = 6.5E-7
+ pkvth0 = 0 stk2 = 0 lodk2 = 1
+ steta0 = 0 lodeta0 = 1

.model nhv_model.4 nmos
+ level = 54 lmin = 1E-6 lmax = 2E-6 wmin = 2E-5
+ wmax = 1.01E-3 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 1.16E-8
+ toxm = 1.16E-8 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 1E23 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {2.1346E-8+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {7.6507E-8-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = -4.1292E-9 dwb = -1.6944E-9 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = 0.778498 lvth0 = 2.005524E-8
+ k1 = 0.88325 k2 = -4.07042E-2 lk2 = 1.305781E-8
+ k3 = -0.884 k3b = 0.43 w0 = 0
+ lpe0 = 2.5E-8 lpeb = -2.182E-7 vbm = -3
+ dvtp0 = 0 dvtp1 = 0 dvt0 = 0
+ dvt1 = 0.53 dvt2 = -0.19251 dvt0w = 0.16
+ dvt1w = 6.9091E6 dvt2w = -0.036016 vfbsdoff = 0
+ u0 = 4.11635E-2 lu0 = 2.637061E-9 ua = -1.424028E-10
+ lua = -7.436395E-18 ub = 1.763188E-18 lub = 1.055951E-25
+ uc = 6.6204E-11 ud = 0 up = 0
+ lp = 1 eu = 1.67 vsat = 1.198856E5
+ lvsat = -2.17495E-2 a0 = 1.702597 la0 = -8.356247E-7
+ ags = 0.152949 lags = 4.284969E-8 b0 = 3.2933E-8
+ b1 = 0 keta = 3.322045E-3 lketa = -2.582464E-8
+ a1 = 0 a2 = 0.659726 rdsw = 724.62
+ rdswmin = 0 rdw = 0 rdwmin = 0
+ rsw = 0 rswmin = 0 prwb = 0.05626
+ prwg = 0.048 wr = 1 voff = -0.20613
+ voffl = -4.257949E-7 minv = 0 nfactor = 0.902098
+ lnfactor = -6.187088E-8 eta0 = 0.032 etab = -0.01932
+ dsub = 0.504 cit = -8E-4 cdsc = 0
+ cdscb = 0 cdscd = 0 pclm = 9.67492E-2
+ lpclm = 2.009904E-7 pdiblc1 = 0.21098 pdiblc2 = 2E-4
+ pdiblcb = -0.26831 drout = 0.36075 pscbe1 = 9.3731E8
+ pscbe2 = 1.68E-6 pvag = 1.99 delta = 0.0246
+ fprout = 10.125 pdits = 0 pditsl = 0
+ pditsd = 0 lambda = 0 vtl = 0
+ lc = 5E-9 xn = 3 alpha0 = 1.4467E-5
+ alpha1 = 0 beta0 = 27.084637 lbeta0 = 4.586737E-6
+ aigbacc = 1 bigbacc = 0 cigbacc = 0
+ nigbacc = 1 aigbinv = 0.35 bigbinv = 0.03
+ cigbinv = 6E-3 eigbinv = 1.1 nigbinv = 3
+ aigc = 0.43 bigc = 0.054 cigc = 0.075
+ aigsd = 0.43 bigsd = 0.054 cigsd = 0.075
+ dlcig = 0 nigc = 1 poxedge = 1
+ pigcd = 1 ntox = 1 toxref = 1.16E-8
+ agidl = 5.06E-11 bgidl = 1.058E9 cgidl = 4E3
+ egidl = 0.8 noia = 2.6E41 noib = 0
+ noic = 0 em = 4.1E7 af = 1
+ ef = 0.89 kf = 0 lintnoi = 0
+ tnoia = 7.5E6 tnoib = 7.2E6 ntnoi = 1
+ rnoia = 0.794 rnoib = 0.38 xpart = 0
+ cgso = {2.754679E-10/sw_func_tox_hv_ratio} cgdo = {2.754679E-10/sw_func_tox_hv_ratio} cgbo = {0/sw_func_tox_hv_ratio}
+ ckappas = 0.6 cf = 0 clc = 1E-7
+ cle = 0.6 dlc = 6.5995E-8 dwc = 0
+ vfbcv = -1 noff = 4 voffcv = -0.4104
+ acde = 0.4176 moin = 15 cgsl = {4.49025E-11/sw_func_tox_hv_ratio}
+ cgdl = {4.49025E-11/sw_func_tox_hv_ratio} ijthsrev = 0.1 ijthsfwd = 0.1
+ xjbvs = 1 bvs = 12.636 jss = 3.75E-4
+ jsws = 5.84E-11 cjs = {8.310E-04*sw_func_nsd_pw_cj} mjs = 0.295
+ mjsws = 0.037586 cjsws = {8.643094E-11*sw_func_nsd_pw_cj} cjswgs = {5.47776E-11*sw_func_nsd_pw_cj}
+ mjswgs = 0.78692 pbs = 0.72468 pbsws = 0.29067
+ pbswgs = 0.54958 xrcrg1 = 12 xrcrg2 = 1
+ rbpb = 50 rbpd = 50 rbps = 50
+ rbdb = 50 rbsb = 50 gbmin = 1E-12
+ tnom = 30 ute = -1.2986 kt1 = -0.3812
+ lkt1 = 1.564371E-8 kt1l = 0 kt2 = -0.019151
+ ua1 = 3.0044E-9 ub1 = -4.006765E-18 lub1 = 4.696243E-25
+ uc1 = -5.9821E-11 at = 9.224112E3 lat = 0.012515
+ prt = 0 njs = 1.0773 xtis = 0.76
+ tpb = 1.344E-3 tpbsw = 9.9005E-4 tpbswg = 0
+ tcj = 6.7434E-4 tcjsw = 2.493E-4 tcjswg = 0
+ tvoff = 0 tvfbsdoff = 0 saref = 3E-6
+ sbref = 3E-6 wlod = 0 ku0 = -4.5E-8
+ kvsat = 0.3 kvth0 = 1.1E-8 tku0 = 0
+ llodku0 = 0 wlodku0 = 1 llodvth = 0
+ wlodvth = 1 lku0 = 0 wku0 = 2E-7
+ pku0 = 0 lkvth0 = 0 wkvth0 = 6.5E-7
+ pkvth0 = 0 stk2 = 0 lodk2 = 1
+ steta0 = 0 lodeta0 = 1

.model nhv_model.5 nmos
+ level = 54 lmin = 8E-7 lmax = 1E-6 wmin = 2E-5
+ wmax = 1.01E-3 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 1.16E-8
+ toxm = 1.16E-8 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 1E23 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {2.1346E-8+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {7.6507E-8-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = -4.1292E-9 dwb = -1.6944E-9 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = 0.788434 lvth0 = 1.163927E-8
+ k1 = 0.88325 k2 = -3.61286E-2 lk2 = 9.182362E-9
+ k3 = -0.884 k3b = 0.43 w0 = 0
+ lpe0 = 2.5E-8 lpeb = -2.182E-7 vbm = -3
+ dvtp0 = 0 dvtp1 = 0 dvt0 = 0
+ dvt1 = 0.53 dvt2 = -0.19251 dvt0w = 0.16
+ dvt1w = 6.9091E6 dvt2w = -0.036016 vfbsdoff = 0
+ u0 = 4.56315E-2 lu0 = -1.147213E-9 ua = -1.607848E-10
+ lua = 8.132965E-18 ub = 1.601827E-18 lub = 2.422655E-25
+ uc = 6.6204E-11 ud = 0 up = 0
+ lp = 1 eu = 1.67 vsat = 8.512623E4
+ lvsat = 7.691287E-3 a0 = -0.597982 la0 = 1.112934E-6
+ ags = 0.34358 lags = -1.18612E-7 b0 = 3.2933E-8
+ b1 = 0 keta = -8.05702E-2 lketa = 4.523094E-8
+ a1 = 0 a2 = 0.659726 rdsw = 724.62
+ rdswmin = 0 rdw = 0 rdwmin = 0
+ rsw = 0 rswmin = 0 prwb = 0.05626
+ prwg = 0.048 wr = 1 voff = -0.20613
+ voffl = -4.257949E-7 minv = 0 nfactor = 0.852374
+ lnfactor = -1.975497E-8 eta0 = 0.032 etab = -0.01932
+ dsub = 0.504 cit = -8E-4 cdsc = 0
+ cdscb = 0 cdscd = 0 pclm = -1.910183
+ lpclm = 1.900834E-6 pdiblc1 = 0.21098 pdiblc2 = 2E-4
+ pdiblcb = -0.26831 drout = 0.36075 pscbe1 = 9.3731E8
+ pscbe2 = 1.68E-6 pvag = 1.99 delta = 0.0246
+ fprout = 10.125 pdits = 0 pditsl = 0
+ pditsd = 0 lambda = 0 vtl = 0
+ lc = 5E-9 xn = 3 alpha0 = 5.108348E-6
+ lalpha0 = 7.926648E-12 alpha1 = 0 beta0 = 22.853439
+ lbeta0 = 8.170502E-6 aigbacc = 1 bigbacc = 0
+ cigbacc = 0 nigbacc = 1 aigbinv = 0.35
+ bigbinv = 0.03 cigbinv = 6E-3 eigbinv = 1.1
+ nigbinv = 3 aigc = 0.43 bigc = 0.054
+ cigc = 0.075 aigsd = 0.43 bigsd = 0.054
+ cigsd = 0.075 dlcig = 0 nigc = 1
+ poxedge = 1 pigcd = 1 ntox = 1
+ toxref = 1.16E-8 agidl = 5.06E-11 bgidl = 1.058E9
+ cgidl = 4E3 egidl = 0.8 noia = 2.6E41
+ noib = 0 noic = 0 em = 4.1E7
+ af = 1 ef = 0.89 kf = 0
+ lintnoi = 0 tnoia = 7.5E6 tnoib = 7.2E6
+ ntnoi = 1 rnoia = 0.794 rnoib = 0.38
+ xpart = 0 cgso = {2.754679E-10/sw_func_tox_hv_ratio} cgdo = {2.754679E-10/sw_func_tox_hv_ratio}
+ cgbo = {0/sw_func_tox_hv_ratio} ckappas = 0.6 cf = 0
+ clc = 1E-7 cle = 0.6 dlc = 6.5995E-8
+ dwc = 0 vfbcv = -1 noff = 4
+ voffcv = -0.4104 acde = 0.4176 moin = 15
+ cgsl = {4.49025E-11/sw_func_tox_hv_ratio} cgdl = {4.49025E-11/sw_func_tox_hv_ratio} ijthsrev = 0.1
+ ijthsfwd = 0.1 xjbvs = 1 bvs = 12.636
+ jss = 3.75E-4 jsws = 5.84E-11 cjs = {8.310E-04*sw_func_nsd_pw_cj}
+ mjs = 0.295 mjsws = 0.037586 cjsws = {8.643094E-11*sw_func_nsd_pw_cj}
+ cjswgs = {5.47776E-11*sw_func_nsd_pw_cj} mjswgs = 0.78692 pbs = 0.72468
+ pbsws = 0.29067 pbswgs = 0.54958 xrcrg1 = 12
+ xrcrg2 = 1 rbpb = 50 rbpd = 50
+ rbps = 50 rbdb = 50 rbsb = 50
+ gbmin = 1E-12 tnom = 30 ute = -1.465199
+ lute = 1.411069E-7 kt1 = -0.336851 lkt1 = -2.191952E-8
+ kt1l = 0 kt2 = -0.019151 ua1 = 6.215715E-9
+ lua1 = -2.719939E-15 ub1 = -9.939305E-18 lub1 = 5.494403E-24
+ uc1 = -5.9821E-11 at = 7.82535E3 lat = 1.36997E-2
+ prt = 0 njs = 1.0773 xtis = 0.76
+ tpb = 1.344E-3 tpbsw = 9.9005E-4 tpbswg = 0
+ tcj = 6.7434E-4 tcjsw = 2.493E-4 tcjswg = 0
+ tvoff = 0 tvfbsdoff = 0 saref = 2.81E-6
+ sbref = 2.81E-6 wlod = 0 ku0 = -4.5E-8
+ kvsat = 0.3 kvth0 = 1.1E-8 tku0 = 0
+ llodku0 = 0 wlodku0 = 1 llodvth = 0
+ wlodvth = 1 lku0 = 0 wku0 = 2E-7
+ pku0 = 0 lkvth0 = 0 wkvth0 = 6.5E-7
+ pkvth0 = 0 stk2 = 0 lodk2 = 1
+ steta0 = 0 lodeta0 = 1

.model nhv_model.6 nmos
+ level = 54 lmin = 6E-7 lmax = 8E-7 wmin = 2E-5
+ wmax = 1.01E-3 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 1.16E-8
+ toxm = 1.16E-8 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 1E23 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {2.1346E-8+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {7.6507E-8-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = -4.1292E-9 dwb = -1.6944E-9 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = 0.806424 k1 = 0.88325
+ k2 = -2.19361E-2 k3 = -0.884 k3b = 0.43
+ w0 = 0 lpe0 = 2.5E-8 lpeb = -2.182E-7
+ vbm = -3 dvtp0 = 0 dvtp1 = 0
+ dvt0 = 0 dvt1 = 0.53 dvt2 = -0.19251
+ dvt0w = 0.16 dvt1w = 6.9091E6 dvt2w = -0.036016
+ vfbsdoff = 0 u0 = 4.38583E-2 ua = -1.482143E-10
+ ub = 1.97628E-18 uc = 6.6204E-11 ud = 0
+ up = 0 lp = 1 eu = 1.67
+ vsat = 9.70141E4 a0 = 1.1222 ags = 0.16025
+ b0 = 3.2933E-8 b1 = 0 keta = -0.01066
+ a1 = 0 a2 = 0.659726 rdsw = 724.62
+ rdswmin = 0 rdw = 0 rdwmin = 0
+ rsw = 0 rswmin = 0 prwb = 0.05626
+ prwg = 0.048 wr = 1 voff = -0.20613
+ voffl = -4.257949E-7 minv = 0 nfactor = 0.82184
+ eta0 = 0.032 etab = -0.01932 dsub = 0.504
+ cit = -8E-4 cdsc = 0 cdscb = 0
+ cdscd = 0 pclm = 1.0278 pdiblc1 = 0.21098
+ pdiblc2 = 2E-4 pdiblcb = -0.26831 drout = 0.36075
+ pscbe1 = 9.3731E8 pscbe2 = 1.68E-6 pvag = 1.99
+ delta = 0.0246 fprout = 10.125 pdits = 0
+ pditsl = 0 pditsd = 0 lambda = 0
+ vtl = 0 lc = 5E-9 xn = 3
+ alpha0 = 1.736E-5 alpha1 = 0 beta0 = 35.482
+ aigbacc = 1 bigbacc = 0 cigbacc = 0
+ nigbacc = 1 aigbinv = 0.35 bigbinv = 0.03
+ cigbinv = 6E-3 eigbinv = 1.1 nigbinv = 3
+ aigc = 0.43 bigc = 0.054 cigc = 0.075
+ aigsd = 0.43 bigsd = 0.054 cigsd = 0.075
+ dlcig = 0 nigc = 1 poxedge = 1
+ pigcd = 1 ntox = 1 toxref = 1.16E-8
+ agidl = 5.06E-11 bgidl = 1.058E9 cgidl = 4E3
+ egidl = 0.8 noia = 2.6E41 noib = 0
+ noic = 0 em = 4.1E7 af = 1
+ ef = 0.89 kf = 0 lintnoi = 0
+ tnoia = 7.5E6 tnoib = 7.2E6 ntnoi = 1
+ rnoia = 0.794 rnoib = 0.38 xpart = 0
+ cgso = {2.754679E-10/sw_func_tox_hv_ratio} cgdo = {2.754679E-10/sw_func_tox_hv_ratio} cgbo = {0/sw_func_tox_hv_ratio}
+ ckappas = 0.6 cf = 0 clc = 1E-7
+ cle = 0.6 dlc = 6.5995E-8 dwc = 0
+ vfbcv = -1 noff = 4 voffcv = -0.4104
+ acde = 0.4176 moin = 15 cgsl = {4.49025E-11/sw_func_tox_hv_ratio}
+ cgdl = {4.49025E-11/sw_func_tox_hv_ratio} ijthsrev = 0.1 ijthsfwd = 0.1
+ xjbvs = 1 bvs = 12.636 jss = 3.75E-4
+ jsws = 5.84E-11 cjs = {8.310E-04*sw_func_nsd_pw_cj} mjs = 0.295
+ mjsws = 0.037586 cjsws = {8.643094E-11*sw_func_nsd_pw_cj} cjswgs = {5.47776E-11*sw_func_nsd_pw_cj}
+ mjswgs = 0.78692 pbs = 0.72468 pbsws = 0.29067
+ pbswgs = 0.54958 xrcrg1 = 12 xrcrg2 = 1
+ rbpb = 50 rbpd = 50 rbps = 50
+ rbdb = 50 rbsb = 50 gbmin = 1E-12
+ tnom = 30 ute = -1.2471 kt1 = -0.37073
+ kt1l = 0 kt2 = -0.019151 ua1 = 2.0117E-9
+ ub1 = -1.447E-18 uc1 = -5.9821E-11 at = 2.9E4
+ prt = 0 njs = 1.0773 xtis = 0.76
+ tpb = 1.344E-3 tpbsw = 9.9005E-4 tpbswg = 0
+ tcj = 6.7434E-4 tcjsw = 2.493E-4 tcjswg = 0
+ tvoff = 0 tvfbsdoff = 0 saref = 2.41E-6
+ sbref = 2.41E-6 wlod = 0 ku0 = -4.5E-8
+ kvsat = 0.3 kvth0 = 1.1E-8 tku0 = 0
+ llodku0 = 0 wlodku0 = 1 llodvth = 0
+ wlodvth = 1 lku0 = 0 wku0 = 2E-7
+ pku0 = 0 lkvth0 = 0 wkvth0 = 6.5E-7
+ pkvth0 = 0 stk2 = 0 lodk2 = 1
+ steta0 = 0 lodeta0 = 1

.model nhv_model.7 nmos
+ level = 54 lmin = 5E-7 lmax = 6E-7 wmin = 2E-5
+ wmax = 1.01E-3 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 1.16E-8
+ toxm = 1.16E-8 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 1E23 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {2.1346E-8+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {7.6507E-8-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = -4.1292E-9 dwb = -1.6944E-9 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = 0.801361 lvth0 = 2.262878E-9
+ k1 = 0.88325 k2 = 2.06956E-2 lk2 = -1.905579E-8
+ k3 = -0.884 k3b = 0.43 w0 = 0
+ lpe0 = 2.5E-8 lpeb = -2.182E-7 vbm = -3
+ dvtp0 = 0 dvtp1 = 0 dvt0 = 0
+ dvt1 = 0.53 dvt2 = -0.19251 dvt0w = 0.16
+ dvt1w = 6.9091E6 dvt2w = -0.036016 vfbsdoff = 0
+ u0 = 2.52481E-2 lu0 = 8.31852E-9 ua = -1.501647E-10
+ lua = 8.718052E-19 ub = -2.513788E-18 lub = 2.006998E-24
+ uc = 6.6204E-11 ud = 0 up = 0
+ lp = 1 eu = 1.67 vsat = 7.509777E4
+ lvsat = 9.796293E-3 a0 = 1.1222 ags = 0.16025
+ b0 = 3.2933E-8 b1 = 0 keta = -0.01066
+ a1 = 0 a2 = 0.659726 rdsw = 724.62
+ rdswmin = 0 rdw = 0 rdwmin = 0
+ rsw = 0 rswmin = 0 prwb = 0.05626
+ prwg = 0.048 wr = 1 voff = -0.20613
+ voffl = -4.257949E-7 minv = 0 nfactor = 1.207411
+ lnfactor = -1.723448E-7 eta0 = 0.032 etab = -0.01932
+ dsub = 0.504 cit = -8E-4 cdsc = 0
+ cdscb = 0 cdscd = 0 pclm = 0.136046
+ lpclm = 3.986016E-7 pdiblc1 = 0.21098 pdiblc2 = 2E-4
+ pdiblcb = -0.26831 drout = 0.36075 pscbe1 = 9.3731E8
+ pscbe2 = 1.68E-6 pvag = 1.99 delta = 0.0246
+ fprout = 10.125 pdits = 0 pditsl = 0
+ pditsd = 0 lambda = 0 vtl = 0
+ lc = 5E-9 xn = 3 alpha0 = 2.73983E-5
+ lalpha0 = -4.486982E-12 alpha1 = 0 beta0 = 30.353547
+ lbeta0 = 2.292347E-6 aigbacc = 1 bigbacc = 0
+ cigbacc = 0 nigbacc = 1 aigbinv = 0.35
+ bigbinv = 0.03 cigbinv = 6E-3 eigbinv = 1.1
+ nigbinv = 3 aigc = 0.43 bigc = 0.054
+ cigc = 0.075 aigsd = 0.43 bigsd = 0.054
+ cigsd = 0.075 dlcig = 0 nigc = 1
+ poxedge = 1 pigcd = 1 ntox = 1
+ toxref = 1.16E-8 agidl = 5.06E-11 bgidl = 1.058E9
+ cgidl = 4E3 egidl = 0.8 noia = 2.6E41
+ noib = 0 noic = 0 em = 4.1E7
+ af = 1 ef = 0.89 kf = 0
+ lintnoi = 0 tnoia = 7.5E6 tnoib = 7.2E6
+ ntnoi = 1 rnoia = 0.794 rnoib = 0.38
+ xpart = 0 cgso = {2.754679E-10/sw_func_tox_hv_ratio} cgdo = {2.754679E-10/sw_func_tox_hv_ratio}
+ cgbo = {0/sw_func_tox_hv_ratio} ckappas = 0.6 cf = 0
+ clc = 1E-7 cle = 0.6 dlc = 6.5995E-8
+ dwc = 0 vfbcv = -1 noff = 4
+ voffcv = -0.4104 acde = 0.4176 moin = 15
+ cgsl = {4.49025E-11/sw_func_tox_hv_ratio} cgdl = {4.49025E-11/sw_func_tox_hv_ratio} ijthsrev = 0.1
+ ijthsfwd = 0.1 xjbvs = 1 bvs = 12.636
+ jss = 3.75E-4 jsws = 5.84E-11 cjs = {8.310E-04*sw_func_nsd_pw_cj}
+ mjs = 0.295 mjsws = 0.037586 cjsws = {8.643094E-11*sw_func_nsd_pw_cj}
+ cjswgs = {5.47776E-11*sw_func_nsd_pw_cj} mjswgs = 0.78692 pbs = 0.72468
+ pbsws = 0.29067 pbswgs = 0.54958 xrcrg1 = 12
+ xrcrg2 = 1 rbpb = 50 rbpd = 50
+ rbps = 50 rbdb = 50 rbsb = 50
+ gbmin = 1E-12 tnom = 30 ute = -1.068402
+ lute = -7.987541E-8 kt1 = -0.440127 lkt1 = 3.101958E-8
+ kt1l = 0 kt2 = -0.019151 ua1 = -1.43283E-9
+ lua1 = 1.539657E-15 ub1 = 5.338311E-18 lub1 = -3.032939E-24
+ uc1 = -5.9821E-11 at = -4.247912E4 lat = 3.19502E-2
+ prt = 0 njs = 1.0773 xtis = 0.76
+ tpb = 1.344E-3 tpbsw = 9.9005E-4 tpbswg = 0
+ tcj = 6.7434E-4 tcjsw = 2.493E-4 tcjswg = 0
+ tvoff = 0 tvfbsdoff = 0 saref = 2.41E-6
+ sbref = 2.41E-6 wlod = 0 ku0 = -4.5E-8
+ kvsat = 0.3 kvth0 = 1.1E-8 tku0 = 0
+ llodku0 = 0 wlodku0 = 1 llodvth = 0
+ wlodvth = 1 lku0 = 0 wku0 = 2E-7
+ pku0 = 0 lkvth0 = 0 wkvth0 = 6.5E-7
+ pkvth0 = 0 stk2 = 0 lodk2 = 1
+ steta0 = 0 lodeta0 = 1

.model nhv_model.8 nmos
+ level = 54 lmin = 8E-6 lmax = 2.02E-5 wmin = 1.5E-5
+ wmax = 2E-5 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 1.16E-8
+ toxm = 1.16E-8 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 1E23 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {2.1346E-8+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {7.6507E-8-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = -4.1292E-9 dwb = -1.6944E-9 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = 0.78882 k1 = 0.88325
+ k2 = -0.039667 k3 = -0.884 k3b = 0.43
+ w0 = 0 lpe0 = 2.5E-8 lpeb = -2.182E-7
+ vbm = -3 dvtp0 = 0 dvtp1 = 0
+ dvt0 = 0 dvt1 = 0.53 dvt2 = -0.19251
+ dvt0w = 0.16 dvt1w = 6.9091E6 dvt2w = -0.036016
+ vfbsdoff = 0 u0 = 4.21082E-2 ua = -5.92431E-11
+ ub = 1.71671E-18 uc = 6.6204E-11 ud = 0
+ up = 0 lp = 1 eu = 1.67
+ vsat = 1.0566E5 a0 = 0.942599 ags = 0.149418
+ b0 = 3.2933E-8 b1 = 0 keta = -0.02132
+ a1 = 0 a2 = 0.659726 rdsw = 724.62
+ rdswmin = 0 rdw = 0 rdwmin = 0
+ rsw = 0 rswmin = 0 prwb = 0.05626
+ prwg = 0.048 wr = 1 voff = -0.20613
+ voffl = -4.257949E-7 minv = 0 nfactor = 0.96538
+ eta0 = 0.032 etab = -0.01932 dsub = 0.504
+ cit = -8E-4 cdsc = 0 cdscb = 0
+ cdscd = 0 pclm = 0.33405 pdiblc1 = 0.21098
+ pdiblc2 = 2E-4 pdiblcb = -0.26831 drout = 0.36075
+ pscbe1 = 9.3731E8 pscbe2 = 1.68E-6 pvag = 1.99
+ delta = 0.0246 fprout = 10.125 pdits = 0
+ pditsl = 0 pditsd = 0 lambda = 0
+ vtl = 0 lc = 5E-9 xn = 3
+ alpha0 = 1.4467E-5 alpha1 = 0 beta0 = 24
+ aigbacc = 1 bigbacc = 0 cigbacc = 0
+ nigbacc = 1 aigbinv = 0.35 bigbinv = 0.03
+ cigbinv = 6E-3 eigbinv = 1.1 nigbinv = 3
+ aigc = 0.43 bigc = 0.054 cigc = 0.075
+ aigsd = 0.43 bigsd = 0.054 cigsd = 0.075
+ dlcig = 0 nigc = 1 poxedge = 1
+ pigcd = 1 ntox = 1 toxref = 1.16E-8
+ agidl = 5.06E-11 bgidl = 1.058E9 cgidl = 4E3
+ egidl = 0.8 noia = 2.6E41 noib = 0
+ noic = 0 em = 4.1E7 af = 1
+ ef = 0.89 kf = 0 lintnoi = 0
+ tnoia = 7.5E6 tnoib = 7.2E6 ntnoi = 1
+ rnoia = 0.794 rnoib = 0.38 xpart = 0
+ cgso = {2.754679E-10/sw_func_tox_hv_ratio} cgdo = {2.754679E-10/sw_func_tox_hv_ratio} cgbo = {0/sw_func_tox_hv_ratio}
+ ckappas = 0.6 cf = 0 clc = 1E-7
+ cle = 0.6 dlc = 6.5995E-8 dwc = 0
+ vfbcv = -1 noff = 4 voffcv = -0.4104
+ acde = 0.4176 moin = 15 cgsl = {4.49025E-11/sw_func_tox_hv_ratio}
+ cgdl = {4.49025E-11/sw_func_tox_hv_ratio} ijthsrev = 0.1 ijthsfwd = 0.1
+ xjbvs = 1 bvs = 12.636 jss = 3.75E-4
+ jsws = 5.84E-11 cjs = {8.310E-04*sw_func_nsd_pw_cj} mjs = 0.295
+ mjsws = 0.037586 cjsws = {8.643094E-11*sw_func_nsd_pw_cj} cjswgs = {5.47776E-11*sw_func_nsd_pw_cj}
+ mjswgs = 0.78692 pbs = 0.72468 pbsws = 0.29067
+ pbswgs = 0.54958 xrcrg1 = 12 xrcrg2 = 1
+ rbpb = 50 rbpd = 50 rbps = 50
+ rbdb = 50 rbsb = 50 gbmin = 1E-12
+ tnom = 30 ute = -1.2986 kt1 = -0.40273
+ kt1l = 0 kt2 = -0.019151 ua1 = 3.0044E-9
+ ub1 = -3.7525E-18 uc1 = -5.9821E-11 at = 1.6E5
+ prt = 0 njs = 1.0773 xtis = 0.76
+ tpb = 1.344E-3 tpbsw = 9.9005E-4 tpbswg = 0
+ tcj = 6.7434E-4 tcjsw = 2.493E-4 tcjswg = 0
+ tvoff = 0 tvfbsdoff = 0 saref = 3E-6
+ sbref = 3E-6 wlod = 0 ku0 = -4.5E-8
+ kvsat = 0.3 kvth0 = 1.1E-8 tku0 = 0
+ llodku0 = 0 wlodku0 = 1 llodvth = 0
+ wlodvth = 1 lku0 = 0 wku0 = 2E-7
+ pku0 = 0 lkvth0 = 0 wkvth0 = 6.5E-7
+ pkvth0 = 0 stk2 = 0 lodk2 = 1
+ steta0 = 0 lodeta0 = 1

.model nhv_model.9 nmos
+ level = 54 lmin = 4E-6 lmax = 8E-6 wmin = 1.5E-5
+ wmax = 2E-5 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 1.16E-8
+ toxm = 1.16E-8 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 1E23 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {2.1346E-8+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {7.6507E-8-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = -4.1292E-9 dwb = -1.6944E-9 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = 0.783367 lvth0 = 4.279042E-8
+ k1 = 0.88325 k2 = -4.10016E-2 lk2 = 1.047271E-8
+ k3 = -0.884 k3b = 0.43 w0 = 0
+ lpe0 = 2.5E-8 lpeb = -2.182E-7 vbm = -3
+ dvtp0 = 0 dvtp1 = 0 dvt0 = 0
+ dvt1 = 0.53 dvt2 = -0.19251 dvt0w = 0.16
+ dvt1w = 6.9091E6 dvt2w = -0.036016 vfbsdoff = 0
+ u0 = 4.15573E-2 lu0 = 4.322814E-9 ua = -1.016037E-10
+ lua = 3.324031E-16 ub = 1.752362E-18 lub = -2.797603E-25
+ uc = 6.6204E-11 ud = 0 up = 0
+ lp = 1 eu = 1.67 vsat = 1.104687E5
+ lvsat = -3.77341E-2 a0 = 1.033611 la0 = -7.141721E-7
+ ags = 0.152066 lags = -2.078241E-8 b0 = 3.2933E-8
+ b1 = 0 keta = -1.72682E-2 lketa = -3.179472E-8
+ a1 = 0 a2 = 0.659726 rdsw = 724.62
+ rdswmin = 0 rdw = 0 rdwmin = 0
+ rsw = 0 rswmin = 0 prwb = 0.05626
+ prwg = 0.048 wr = 1 voff = -0.20613
+ voffl = -4.257949E-7 minv = 0 nfactor = 1.012092
+ lnfactor = -3.665486E-7 eta0 = 0.032 etab = -0.01932
+ dsub = 0.504 cit = -8E-4 cdsc = 0
+ cdscb = 0 cdscd = 0 pclm = 0.259909
+ lpclm = 5.817837E-7 pdiblc1 = 0.21098 pdiblc2 = 2E-4
+ pdiblcb = -0.26831 drout = 0.36075 pscbe1 = 9.3731E8
+ pscbe2 = 1.68E-6 pvag = 1.99 delta = 0.0246
+ fprout = 10.125 pdits = 0 pditsl = 0
+ pditsd = 0 lambda = 0 vtl = 0
+ lc = 5E-9 xn = 3 alpha0 = 1.4467E-5
+ alpha1 = 0 beta0 = 21.499459 lbeta0 = 1.962171E-5
+ aigbacc = 1 bigbacc = 0 cigbacc = 0
+ nigbacc = 1 aigbinv = 0.35 bigbinv = 0.03
+ cigbinv = 6E-3 eigbinv = 1.1 nigbinv = 3
+ aigc = 0.43 bigc = 0.054 cigc = 0.075
+ aigsd = 0.43 bigsd = 0.054 cigsd = 0.075
+ dlcig = 0 nigc = 1 poxedge = 1
+ pigcd = 1 ntox = 1 toxref = 1.16E-8
+ agidl = 5.06E-11 bgidl = 1.058E9 cgidl = 4E3
+ egidl = 0.8 noia = 2.6E41 noib = 0
+ noic = 0 em = 4.1E7 af = 1
+ ef = 0.89 kf = 0 lintnoi = 0
+ tnoia = 7.5E6 tnoib = 7.2E6 ntnoi = 1
+ rnoia = 0.794 rnoib = 0.38 xpart = 0
+ cgso = {2.754679E-10/sw_func_tox_hv_ratio} cgdo = {2.754679E-10/sw_func_tox_hv_ratio} cgbo = {0/sw_func_tox_hv_ratio}
+ ckappas = 0.6 cf = 0 clc = 1E-7
+ cle = 0.6 dlc = 6.5995E-8 dwc = 0
+ vfbcv = -1 noff = 4 voffcv = -0.4104
+ acde = 0.4176 moin = 15 cgsl = {4.49025E-11/sw_func_tox_hv_ratio}
+ cgdl = {4.49025E-11/sw_func_tox_hv_ratio} ijthsrev = 0.1 ijthsfwd = 0.1
+ xjbvs = 1 bvs = 12.636 jss = 3.75E-4
+ jsws = 5.84E-11 cjs = {8.310E-04*sw_func_nsd_pw_cj} mjs = 0.295
+ mjsws = 0.037586 cjsws = {8.643094E-11*sw_func_nsd_pw_cj} cjswgs = {5.47776E-11*sw_func_nsd_pw_cj}
+ mjswgs = 0.78692 pbs = 0.72468 pbsws = 0.29067
+ pbswgs = 0.54958 xrcrg1 = 12 xrcrg2 = 1
+ rbpb = 50 rbpd = 50 rbps = 50
+ rbdb = 50 rbsb = 50 gbmin = 1E-12
+ tnom = 30 ute = -1.33707 lute = 3.018725E-7
+ kt1 = -0.414271 lkt1 = 9.056174E-8 kt1l = 0
+ kt2 = -0.019151 ua1 = 3.0044E-9 ub1 = -3.7525E-18
+ uc1 = -5.9821E-11 at = 2.369397E5 lat = -0.603745
+ prt = 0 njs = 1.0773 xtis = 0.76
+ tpb = 1.344E-3 tpbsw = 9.9005E-4 tpbswg = 0
+ tcj = 6.7434E-4 tcjsw = 2.493E-4 tcjswg = 0
+ tvoff = 0 tvfbsdoff = 0 saref = 3E-6
+ sbref = 3E-6 wlod = 0 ku0 = -4.5E-8
+ kvsat = 0.3 kvth0 = 1.1E-8 tku0 = 0
+ llodku0 = 0 wlodku0 = 1 llodvth = 0
+ wlodvth = 1 lku0 = 0 wku0 = 2E-7
+ pku0 = 0 lkvth0 = 0 wkvth0 = 6.5E-7
+ pkvth0 = 0 stk2 = 0 lodk2 = 1
+ steta0 = 0 lodeta0 = 1

.model nhv_model.10 nmos
+ level = 54 lmin = 2E-6 lmax = 4E-6 wmin = 1.5E-5
+ wmax = 2E-5 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 1.16E-8
+ toxm = 1.16E-8 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 1E23 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {2.1346E-8+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {7.6507E-8-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = -4.1292E-9 dwb = -1.6944E-9 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = 0.799231 lvth0 = -1.823938E-8
+ k1 = 0.88325 k2 = -4.25688E-2 lk2 = 1.650177E-8
+ k3 = -0.884 k3b = 0.43 w0 = 0
+ lpe0 = 2.5E-8 lpeb = -2.182E-7 vbm = -3
+ dvtp0 = 0 dvtp1 = 0 dvt0 = 0
+ dvt1 = 0.53 dvt2 = -0.19251 dvt0w = 0.16
+ dvt1w = 6.9091E6 dvt2w = -0.036016 vfbsdoff = 0
+ u0 = 4.27638E-2 lu0 = -3.18674E-10 ua = 1.059937E-10
+ lua = -4.662212E-16 ub = 1.549686E-18 lub = 4.99931E-25
+ uc = 6.6204E-11 ud = 0 up = 0
+ lp = 1 eu = 1.67 vsat = 9.377998E4
+ lvsat = 2.64674E-2 a0 = 0.476534 la0 = 1.428898E-6
+ ags = 0.119435 lags = 1.047503E-7 b0 = 3.2933E-8
+ b1 = 0 keta = -3.92681E-2 lketa = 5.283878E-8
+ a1 = 0 a2 = 0.659726 rdsw = 724.62
+ rdswmin = 0 rdw = 0 rdwmin = 0
+ rsw = 0 rswmin = 0 prwb = 0.05626
+ prwg = 0.048 wr = 1 voff = -0.20613
+ voffl = -4.257949E-7 minv = 0 nfactor = 0.961332
+ lnfactor = -1.71274E-7 eta0 = 0.032 etab = -0.01932
+ dsub = 0.504 cit = -8E-4 cdsc = 0
+ cdscb = 0 cdscd = 0 pclm = 0.600982
+ lpclm = -7.303213E-7 pdiblc1 = 0.21098 pdiblc2 = 2E-4
+ pdiblcb = -0.26831 drout = 0.36075 pscbe1 = 9.3731E8
+ pscbe2 = 1.68E-6 pvag = 1.99 delta = 0.0246
+ fprout = 10.125 pdits = 0 pditsl = 0
+ pditsd = 0 lambda = 0 vtl = 0
+ lc = 5E-9 xn = 3 alpha0 = 1.4467E-5
+ alpha1 = 0 beta0 = 23.859073 lbeta0 = 1.054431E-5
+ aigbacc = 1 bigbacc = 0 cigbacc = 0
+ nigbacc = 1 aigbinv = 0.35 bigbinv = 0.03
+ cigbinv = 6E-3 eigbinv = 1.1 nigbinv = 3
+ aigc = 0.43 bigc = 0.054 cigc = 0.075
+ aigsd = 0.43 bigsd = 0.054 cigsd = 0.075
+ dlcig = 0 nigc = 1 poxedge = 1
+ pigcd = 1 ntox = 1 toxref = 1.16E-8
+ agidl = 5.06E-11 bgidl = 1.058E9 cgidl = 4E3
+ egidl = 0.8 noia = 2.6E41 noib = 0
+ noic = 0 em = 4.1E7 af = 1
+ ef = 0.89 kf = 0 lintnoi = 0
+ tnoia = 7.5E6 tnoib = 7.2E6 ntnoi = 1
+ rnoia = 0.794 rnoib = 0.38 xpart = 0
+ cgso = {2.754679E-10/sw_func_tox_hv_ratio} cgdo = {2.754679E-10/sw_func_tox_hv_ratio} cgbo = {0/sw_func_tox_hv_ratio}
+ ckappas = 0.6 cf = 0 clc = 1E-7
+ cle = 0.6 dlc = 6.5995E-8 dwc = 0
+ vfbcv = -1 noff = 4 voffcv = -0.4104
+ acde = 0.4176 moin = 15 cgsl = {4.49025E-11/sw_func_tox_hv_ratio}
+ cgdl = {4.49025E-11/sw_func_tox_hv_ratio} ijthsrev = 0.1 ijthsfwd = 0.1
+ xjbvs = 1 bvs = 12.636 jss = 3.75E-4
+ jsws = 5.84E-11 cjs = {8.310E-04*sw_func_nsd_pw_cj} mjs = 0.295
+ mjsws = 0.037586 cjsws = {8.643094E-11*sw_func_nsd_pw_cj} cjswgs = {5.47776E-11*sw_func_nsd_pw_cj}
+ mjswgs = 0.78692 pbs = 0.72468 pbsws = 0.29067
+ pbswgs = 0.54958 xrcrg1 = 12 xrcrg2 = 1
+ rbpb = 50 rbpd = 50 rbps = 50
+ rbdb = 50 rbsb = 50 gbmin = 1E-12
+ tnom = 30 ute = -1.22166 lute = -1.421066E-7
+ kt1 = -0.407353 lkt1 = 6.394796E-8 kt1l = 0
+ kt2 = -0.019151 ua1 = 3.0044E-9 ub1 = -3.7525E-18
+ uc1 = -5.9821E-11 at = 1.391036E5 lat = -0.227371
+ prt = 0 njs = 1.0773 xtis = 0.76
+ tpb = 1.344E-3 tpbsw = 9.9005E-4 tpbswg = 0
+ tcj = 6.7434E-4 tcjsw = 2.493E-4 tcjswg = 0
+ tvoff = 0 tvfbsdoff = 0 saref = 3E-6
+ sbref = 3E-6 wlod = 0 ku0 = -4.5E-8
+ kvsat = 0.3 kvth0 = 1.1E-8 tku0 = 0
+ llodku0 = 0 wlodku0 = 1 llodvth = 0
+ wlodvth = 1 lku0 = 0 wku0 = 2E-7
+ pku0 = 0 lkvth0 = 0 wkvth0 = 6.5E-7
+ pkvth0 = 0 stk2 = 0 lodk2 = 1
+ steta0 = 0 lodeta0 = 1

.model nhv_model.11 nmos
+ level = 54 lmin = 1E-6 lmax = 2E-6 wmin = 1.5E-5
+ wmax = 2E-5 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 1.16E-8
+ toxm = 1.16E-8 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 1E23 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {2.1346E-8+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {7.6507E-8-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = -4.1292E-9 dwb = -1.6944E-9 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = 0.779602 lvth0 = 1.801487E-8
+ wvth0 = -2.204693E-8 pvth0 = 4.072037E-14 k1 = 0.88325
+ k2 = -4.00796E-2 lk2 = 1.190425E-8 wk2 = -1.246461E-8
+ pk2 = 2.302195E-14 k3 = -0.884 k3b = 0.43
+ w0 = 0 lpe0 = 2.5E-8 lpeb = -2.182E-7
+ vbm = -3 dvtp0 = 0 dvtp1 = 0
+ dvt0 = 0 dvt1 = 0.53 dvt2 = -0.19251
+ dvt0w = 0.16 dvt1w = 6.9091E6 dvt2w = -0.036016
+ vfbsdoff = 0 u0 = 4.05272E-2 lu0 = 3.812428E-9
+ wu0 = 1.270024E-8 pu0 = -2.345717E-14 ua = -1.49239E-10
+ lua = 5.190056E-18 wua = 1.364331E-16 pua = -2.5199E-22
+ ub = 1.659382E-18 lub = 2.973247E-25 wub = 2.071703E-24
+ pub = -3.826407E-30 uc = 6.6204E-11 ud = 0
+ up = 0 lp = 1 eu = 1.67
+ vsat = 1.274868E5 lvsat = -3.57887E-2 wvsat = -0.151699
+ pvsat = 2.80186E-7 a0 = 1.759572 la0 = -9.408556E-7
+ wa0 = -1.137055E-6 pa0 = 2.100125E-12 ags = 3.84106E-2
+ lags = 2.544009E-7 wags = 2.285882E-6 pags = -4.221993E-12
+ b0 = 3.2933E-8 b1 = 0 keta = 3.322045E-3
+ lketa = -2.582464E-8 a1 = 0 a2 = 0.659726
+ rdsw = 724.62 rdswmin = 0 rdw = 0
+ rdwmin = 0 rsw = 0 rswmin = 0
+ prwb = 0.05626 prwg = 0.048 wr = 1
+ voff = -0.20613 voffl = -4.257949E-7 minv = 0
+ nfactor = 0.90334 lnfactor = -6.416397E-8 wnfactor = -2.477751E-8
+ pnfactor = 4.576372E-14 eta0 = 0.032 etab = -0.01932
+ dsub = 0.504 cit = -8E-4 cdsc = 0
+ cdscb = 0 cdscd = 0 pclm = 9.67492E-2
+ lpclm = 2.009904E-7 pdiblc1 = 0.21098 pdiblc2 = 2E-4
+ pdiblcb = -0.26831 drout = 0.36075 pscbe1 = 9.3731E8
+ pscbe2 = 1.68E-6 pvag = 1.99 delta = 0.0246
+ fprout = 10.125 pdits = 0 pditsl = 0
+ pditsd = 0 lambda = 0 vtl = 0
+ lc = 5E-9 xn = 3 alpha0 = 1.4467E-5
+ alpha1 = 0 beta0 = 27.14798 lbeta0 = 4.469743E-6
+ wbeta0 = -1.264159E-6 pbeta0 = 2.334884E-12 aigbacc = 1
+ bigbacc = 0 cigbacc = 0 nigbacc = 1
+ aigbinv = 0.35 bigbinv = 0.03 cigbinv = 6E-3
+ eigbinv = 1.1 nigbinv = 3 aigc = 0.43
+ bigc = 0.054 cigc = 0.075 aigsd = 0.43
+ bigsd = 0.054 cigsd = 0.075 dlcig = 0
+ nigc = 1 poxedge = 1 pigcd = 1
+ ntox = 1 toxref = 1.16E-8 agidl = 5.06E-11
+ bgidl = 1.058E9 cgidl = 4E3 egidl = 0.8
+ noia = 2.6E41 noib = 0 noic = 0
+ em = 4.1E7 af = 1 ef = 0.89
+ kf = 0 lintnoi = 0 tnoia = 7.5E6
+ tnoib = 7.2E6 ntnoi = 1 rnoia = 0.794
+ rnoib = 0.38 xpart = 0 cgso = {2.754679E-10/sw_func_tox_hv_ratio}
+ cgdo = {2.754679E-10/sw_func_tox_hv_ratio} cgbo = {0/sw_func_tox_hv_ratio} ckappas = 0.6
+ cf = 0 clc = 1E-7 cle = 0.6
+ dlc = 6.5995E-8 dwc = 0 vfbcv = -1
+ noff = 4 voffcv = -0.4104 acde = 0.4176
+ moin = 15 cgsl = {4.49025E-11/sw_func_tox_hv_ratio} cgdl = {4.49025E-11/sw_func_tox_hv_ratio}
+ ijthsrev = 0.1 ijthsfwd = 0.1 xjbvs = 1
+ bvs = 12.636 jss = 3.75E-4 jsws = 5.84E-11
+ cjs = {8.310E-04*sw_func_nsd_pw_cj} mjs = 0.295 mjsws = 0.037586
+ cjsws = {8.643094E-11*sw_func_nsd_pw_cj} cjswgs = {5.47776E-11*sw_func_nsd_pw_cj} mjswgs = 0.78692
+ pbs = 0.72468 pbsws = 0.29067 pbswgs = 0.54958
+ xrcrg1 = 12 xrcrg2 = 1 rbpb = 50
+ rbpd = 50 rbps = 50 rbdb = 50
+ rbsb = 50 gbmin = 1E-12 tnom = 30
+ ute = -1.2986 kt1 = -0.3812 lkt1 = 1.564371E-8
+ kt1l = 0 kt2 = -0.019151 ua1 = 3.0044E-9
+ ub1 = -4.006765E-18 lub1 = 4.696243E-25 uc1 = -5.9821E-11
+ at = 9.224112E3 lat = 0.012515 prt = 0
+ njs = 1.0773 xtis = 0.76 tpb = 1.344E-3
+ tpbsw = 9.9005E-4 tpbswg = 0 tcj = 6.7434E-4
+ tcjsw = 2.493E-4 tcjswg = 0 tvoff = 0
+ tvfbsdoff = 0 saref = 3E-6 sbref = 3E-6
+ wlod = 0 ku0 = -4.5E-8 kvsat = 0.3
+ kvth0 = 1.1E-8 tku0 = 0 llodku0 = 0
+ wlodku0 = 1 llodvth = 0 wlodvth = 1
+ lku0 = 0 wku0 = 2E-7 pku0 = 0
+ lkvth0 = 0 wkvth0 = 6.5E-7 pkvth0 = 0
+ stk2 = 0 lodk2 = 1 steta0 = 0
+ lodeta0 = 1

.model nhv_model.12 nmos
+ level = 54 lmin = 8E-7 lmax = 1E-6 wmin = 1.5E-5
+ wmax = 2E-5 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 1.16E-8
+ toxm = 1.16E-8 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 1E23 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {2.1346E-8+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {7.6507E-8-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = -4.1292E-9 dwb = -1.6944E-9 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = 0.78291 lvth0 = 1.521291E-8
+ wvth0 = 1.102346E-7 pvth0 = -7.132027E-14 k1 = 0.88325
+ k2 = -3.92514E-2 lk2 = 1.120278E-8 wk2 = 6.232303E-8
+ pk2 = -4.032213E-14 k3 = -0.884 k3b = 0.43
+ w0 = 0 lpe0 = 2.5E-8 lpeb = -2.182E-7
+ vbm = -3 dvtp0 = 0 dvtp1 = 0
+ dvt0 = 0 dvt1 = 0.53 dvt2 = -0.19251
+ dvt0w = 0.16 dvt1w = 6.9091E6 dvt2w = -0.036016
+ vfbsdoff = 0 u0 = 4.88133E-2 lu0 = -3.205828E-9
+ wu0 = -6.350122E-8 pu0 = 4.10844E-14 ua = -1.266036E-10
+ lua = -1.398181E-17 wua = -6.821654E-16 pua = 4.413514E-22
+ ub = 2.120861E-18 lub = -9.354206E-26 wub = -1.035852E-23
+ pub = 6.701816E-30 uc = 6.6204E-11 ud = 0
+ up = 0 lp = 1 eu = 1.67
+ vsat = 4.712034E4 lvsat = 3.22806E-2 wvsat = 0.758495
+ pvsat = -4.907358E-7 a0 = -0.882854 la0 = 1.297242E-6
+ wa0 = 5.685276E-6 pa0 = -3.678294E-12 ags = 0.916273
+ lags = -4.891364E-7 wags = -1.142941E-5 pags = 7.394669E-12
+ b0 = 3.2933E-8 b1 = 0 keta = -8.05702E-2
+ lketa = 4.523094E-8 a1 = 0 a2 = 0.659726
+ rdsw = 724.62 rdswmin = 0 rdw = 0
+ rdwmin = 0 rsw = 0 rswmin = 0
+ prwb = 0.05626 prwg = 0.048 wr = 1
+ voff = -0.20613 voffl = -4.257949E-7 minv = 0
+ nfactor = 0.846166 lnfactor = -1.573872E-8 wnfactor = 1.238876E-7
+ pnfactor = -8.015352E-14 eta0 = 0.032 etab = -0.01932
+ dsub = 0.504 cit = -8E-4 cdsc = 0
+ cdscb = 0 cdscd = 0 pclm = -1.910183
+ lpclm = 1.900834E-6 pdiblc1 = 0.21098 pdiblc2 = 2E-4
+ pdiblcb = -0.26831 drout = 0.36075 pscbe1 = 9.3731E8
+ pscbe2 = 1.68E-6 pvag = 1.99 delta = 0.0246
+ fprout = 10.125 pdits = 0 pditsl = 0
+ pditsd = 0 lambda = 0 vtl = 0
+ lc = 5E-9 xn = 3 alpha0 = 5.108348E-6
+ lalpha0 = 7.926648E-12 alpha1 = 0 beta0 = 22.536723
+ lbeta0 = 8.375413E-6 wbeta0 = 6.320794E-6 pbeta0 = -4.089465E-12
+ aigbacc = 1 bigbacc = 0 cigbacc = 0
+ nigbacc = 1 aigbinv = 0.35 bigbinv = 0.03
+ cigbinv = 6E-3 eigbinv = 1.1 nigbinv = 3
+ aigc = 0.43 bigc = 0.054 cigc = 0.075
+ aigsd = 0.43 bigsd = 0.054 cigsd = 0.075
+ dlcig = 0 nigc = 1 poxedge = 1
+ pigcd = 1 ntox = 1 toxref = 1.16E-8
+ agidl = 5.06E-11 bgidl = 1.058E9 cgidl = 4E3
+ egidl = 0.8 noia = 2.6E41 noib = 0
+ noic = 0 em = 4.1E7 af = 1
+ ef = 0.89 kf = 0 lintnoi = 0
+ tnoia = 7.5E6 tnoib = 7.2E6 ntnoi = 1
+ rnoia = 0.794 rnoib = 0.38 xpart = 0
+ cgso = {2.754679E-10/sw_func_tox_hv_ratio} cgdo = {2.754679E-10/sw_func_tox_hv_ratio} cgbo = {0/sw_func_tox_hv_ratio}
+ ckappas = 0.6 cf = 0 clc = 1E-7
+ cle = 0.6 dlc = 6.5995E-8 dwc = 0
+ vfbcv = -1 noff = 4 voffcv = -0.4104
+ acde = 0.4176 moin = 15 cgsl = {4.49025E-11/sw_func_tox_hv_ratio}
+ cgdl = {4.49025E-11/sw_func_tox_hv_ratio} ijthsrev = 0.1 ijthsfwd = 0.1
+ xjbvs = 1 bvs = 12.636 jss = 3.75E-4
+ jsws = 5.84E-11 cjs = {8.310E-04*sw_func_nsd_pw_cj} mjs = 0.295
+ mjsws = 0.037586 cjsws = {8.643094E-11*sw_func_nsd_pw_cj} cjswgs = {5.47776E-11*sw_func_nsd_pw_cj}
+ mjswgs = 0.78692 pbs = 0.72468 pbsws = 0.29067
+ pbswgs = 0.54958 xrcrg1 = 12 xrcrg2 = 1
+ rbpb = 50 rbpd = 50 rbps = 50
+ rbdb = 50 rbsb = 50 gbmin = 1E-12
+ tnom = 30 ute = -1.465199 lute = 1.411069E-7
+ kt1 = -0.336851 lkt1 = -2.191952E-8 kt1l = 0
+ kt2 = -0.019151 ua1 = 6.215715E-9 lua1 = -2.719939E-15
+ ub1 = -9.939305E-18 lub1 = 5.494403E-24 uc1 = -5.9821E-11
+ at = 7.82535E3 lat = 1.36997E-2 prt = 0
+ njs = 1.0773 xtis = 0.76 tpb = 1.344E-3
+ tpbsw = 9.9005E-4 tpbswg = 0 tcj = 6.7434E-4
+ tcjsw = 2.493E-4 tcjswg = 0 tvoff = 0
+ tvfbsdoff = 0 saref = 2.81E-6 sbref = 2.81E-6
+ wlod = 0 ku0 = -4.5E-8 kvsat = 0.3
+ kvth0 = 1.1E-8 tku0 = 0 llodku0 = 0
+ wlodku0 = 1 llodvth = 0 wlodvth = 1
+ lku0 = 0 wku0 = 2E-7 pku0 = 0
+ lkvth0 = 0 wkvth0 = 6.5E-7 pkvth0 = 0
+ stk2 = 0 lodk2 = 1 steta0 = 0
+ lodeta0 = 1

.model nhv_model.13 nmos
+ level = 54 lmin = 6E-7 lmax = 8E-7 wmin = 1.5E-5
+ wmax = 2E-5 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 1.16E-8
+ toxm = 1.16E-8 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 1E23 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {2.1346E-8+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {7.6507E-8-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = -4.1292E-9 dwb = -1.6944E-9 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = 0.806424 k1 = 0.88325
+ k2 = -2.19361E-2 k3 = -0.884 k3b = 0.43
+ w0 = 0 lpe0 = 2.5E-8 lpeb = -2.182E-7
+ vbm = -3 dvtp0 = 0 dvtp1 = 0
+ dvt0 = 0 dvt1 = 0.53 dvt2 = -0.19251
+ dvt0w = 0.16 dvt1w = 6.9091E6 dvt2w = -0.036016
+ vfbsdoff = 0 u0 = 4.38583E-2 ua = -1.482143E-10
+ ub = 1.97628E-18 uc = 6.6204E-11 ud = 0
+ up = 0 lp = 1 eu = 1.67
+ vsat = 9.70141E4 a0 = 1.1222 ags = 0.16025
+ b0 = 3.2933E-8 b1 = 0 keta = -0.01066
+ a1 = 0 a2 = 0.659726 rdsw = 724.62
+ rdswmin = 0 rdw = 0 rdwmin = 0
+ rsw = 0 rswmin = 0 prwb = 0.05626
+ prwg = 0.048 wr = 1 voff = -0.20613
+ voffl = -4.257949E-7 minv = 0 nfactor = 0.82184
+ eta0 = 0.032 etab = -0.01932 dsub = 0.504
+ cit = -8E-4 cdsc = 0 cdscb = 0
+ cdscd = 0 pclm = 1.0278 pdiblc1 = 0.21098
+ pdiblc2 = 2E-4 pdiblcb = -0.26831 drout = 0.36075
+ pscbe1 = 9.3731E8 pscbe2 = 1.68E-6 pvag = 1.99
+ delta = 0.0246 fprout = 10.125 pdits = 0
+ pditsl = 0 pditsd = 0 lambda = 0
+ vtl = 0 lc = 5E-9 xn = 3
+ alpha0 = 1.736E-5 alpha1 = 0 beta0 = 35.482
+ aigbacc = 1 bigbacc = 0 cigbacc = 0
+ nigbacc = 1 aigbinv = 0.35 bigbinv = 0.03
+ cigbinv = 6E-3 eigbinv = 1.1 nigbinv = 3
+ aigc = 0.43 bigc = 0.054 cigc = 0.075
+ aigsd = 0.43 bigsd = 0.054 cigsd = 0.075
+ dlcig = 0 nigc = 1 poxedge = 1
+ pigcd = 1 ntox = 1 toxref = 1.16E-8
+ agidl = 5.06E-11 bgidl = 1.058E9 cgidl = 4E3
+ egidl = 0.8 noia = 2.6E41 noib = 0
+ noic = 0 em = 4.1E7 af = 1
+ ef = 0.89 kf = 0 lintnoi = 0
+ tnoia = 7.5E6 tnoib = 7.2E6 ntnoi = 1
+ rnoia = 0.794 rnoib = 0.38 xpart = 0
+ cgso = {2.754679E-10/sw_func_tox_hv_ratio} cgdo = {2.754679E-10/sw_func_tox_hv_ratio} cgbo = {0/sw_func_tox_hv_ratio}
+ ckappas = 0.6 cf = 0 clc = 1E-7
+ cle = 0.6 dlc = 6.5995E-8 dwc = 0
+ vfbcv = -1 noff = 4 voffcv = -0.4104
+ acde = 0.4176 moin = 15 cgsl = {4.49025E-11/sw_func_tox_hv_ratio}
+ cgdl = {4.49025E-11/sw_func_tox_hv_ratio} ijthsrev = 0.1 ijthsfwd = 0.1
+ xjbvs = 1 bvs = 12.636 jss = 3.75E-4
+ jsws = 5.84E-11 cjs = {8.310E-04*sw_func_nsd_pw_cj} mjs = 0.295
+ mjsws = 0.037586 cjsws = {8.643094E-11*sw_func_nsd_pw_cj} cjswgs = {5.47776E-11*sw_func_nsd_pw_cj}
+ mjswgs = 0.78692 pbs = 0.72468 pbsws = 0.29067
+ pbswgs = 0.54958 xrcrg1 = 12 xrcrg2 = 1
+ rbpb = 50 rbpd = 50 rbps = 50
+ rbdb = 50 rbsb = 50 gbmin = 1E-12
+ tnom = 30 ute = -1.2471 kt1 = -0.37073
+ kt1l = 0 kt2 = -0.019151 ua1 = 2.0117E-9
+ ub1 = -1.447E-18 uc1 = -5.9821E-11 at = 2.9E4
+ prt = 0 njs = 1.0773 xtis = 0.76
+ tpb = 1.344E-3 tpbsw = 9.9005E-4 tpbswg = 0
+ tcj = 6.7434E-4 tcjsw = 2.493E-4 tcjswg = 0
+ tvoff = 0 tvfbsdoff = 0 saref = 2.41E-6
+ sbref = 2.41E-6 wlod = 0 ku0 = -4.5E-8
+ kvsat = 0.3 kvth0 = 1.1E-8 tku0 = 0
+ llodku0 = 0 wlodku0 = 1 llodvth = 0
+ wlodvth = 1 lku0 = 0 wku0 = 2E-7
+ pku0 = 0 lkvth0 = 0 wkvth0 = 6.5E-7
+ pkvth0 = 0 stk2 = 0 lodk2 = 1
+ steta0 = 0 lodeta0 = 1

.model nhv_model.14 nmos
+ level = 54 lmin = 5E-7 lmax = 6E-7 wmin = 1.5E-5
+ wmax = 2E-5 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 1.16E-8
+ toxm = 1.16E-8 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 1E23 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {2.1346E-8+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {7.6507E-8-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = -4.1292E-9 dwb = -1.6944E-9 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = 0.834006 lvth0 = -1.232896E-8
+ wvth0 = -6.515054E-7 pvth0 = 2.912138E-13 k1 = 0.88325
+ k2 = 2.50801E-2 lk2 = -2.10156E-8 wk2 = -8.750266E-8
+ pk2 = 3.911246E-14 k3 = -0.884 k3b = 0.43
+ w0 = 0 lpe0 = 2.5E-8 lpeb = -2.182E-7
+ vbm = -3 dvtp0 = 0 dvtp1 = 0
+ dvt0 = 0 dvt1 = 0.53 dvt2 = -0.19251
+ dvt0w = 0.16 dvt1w = 6.9091E6 dvt2w = -0.036016
+ vfbsdoff = 0 u0 = 0.030821 lu0 = 5.827468E-9
+ wu0 = -1.11222E-7 pu0 = 4.971468E-14 ua = -2.076167E-10
+ lua = 2.655205E-17 wua = 1.146587E-15 pua = -5.125085E-22
+ ub = -4.561857E-18 lub = 2.922456E-24 wub = 4.087393E-23
+ pub = -1.827008E-29 uc = 6.6204E-11 ud = 0
+ up = 0 lp = 1 eu = 1.67
+ vsat = 9.678782E4 lvsat = 1.011423E-4 wvsat = -0.432875
+ pvsat = 1.934891E-7 a0 = 1.1222 ags = 0.16025
+ b0 = 3.2933E-8 b1 = 0 keta = -0.01066
+ a1 = 0 a2 = 0.659726 rdsw = 724.62
+ rdswmin = 0 rdw = 0 rdwmin = 0
+ rsw = 0 rswmin = 0 prwb = 0.05626
+ prwg = 0.048 wr = 1 voff = -0.20613
+ voffl = -4.257949E-7 minv = 0 nfactor = 1.511959
+ lnfactor = -3.084734E-7 wnfactor = -6.077955E-6 pnfactor = 2.716761E-12
+ eta0 = 0.032 etab = -0.01932 dsub = 0.504
+ cit = -8E-4 cdsc = 0 cdscb = 0
+ cdscd = 0 pclm = -1.998072 lpclm = 1.352523E-6
+ wpclm = 4.259126E-5 ppclm = -1.90377E-11 pdiblc1 = 0.21098
+ pdiblc2 = 2E-4 pdiblcb = -0.26831 drout = 0.36075
+ pscbe1 = 9.3731E8 pscbe2 = 1.68E-6 pvag = 1.99
+ delta = 0.0246 fprout = 10.125 pdits = 0
+ pditsl = 0 pditsd = 0 lambda = 0
+ vtl = 0 lc = 5E-9 xn = 3
+ alpha0 = 2.73983E-5 lalpha0 = -4.486982E-12 alpha1 = 0
+ beta0 = 30.353547 lbeta0 = 2.292347E-6 aigbacc = 1
+ bigbacc = 0 cigbacc = 0 nigbacc = 1
+ aigbinv = 0.35 bigbinv = 0.03 cigbinv = 6E-3
+ eigbinv = 1.1 nigbinv = 3 aigc = 0.43
+ bigc = 0.054 cigc = 0.075 aigsd = 0.43
+ bigsd = 0.054 cigsd = 0.075 dlcig = 0
+ nigc = 1 poxedge = 1 pigcd = 1
+ ntox = 1 toxref = 1.16E-8 agidl = 5.06E-11
+ bgidl = 1.058E9 cgidl = 4E3 egidl = 0.8
+ noia = 2.6E41 noib = 0 noic = 0
+ em = 4.1E7 af = 1 ef = 0.89
+ kf = 0 lintnoi = 0 tnoia = 7.5E6
+ tnoib = 7.2E6 ntnoi = 1 rnoia = 0.794
+ rnoib = 0.38 xpart = 0 cgso = {2.754679E-10/sw_func_tox_hv_ratio}
+ cgdo = {2.754679E-10/sw_func_tox_hv_ratio} cgbo = {0/sw_func_tox_hv_ratio} ckappas = 0.6
+ cf = 0 clc = 1E-7 cle = 0.6
+ dlc = 6.5995E-8 dwc = 0 vfbcv = -1
+ noff = 4 voffcv = -0.4104 acde = 0.4176
+ moin = 15 cgsl = {4.49025E-11/sw_func_tox_hv_ratio} cgdl = {4.49025E-11/sw_func_tox_hv_ratio}
+ ijthsrev = 0.1 ijthsfwd = 0.1 xjbvs = 1
+ bvs = 12.636 jss = 3.75E-4 jsws = 5.84E-11
+ cjs = {8.310E-04*sw_func_nsd_pw_cj} mjs = 0.295 mjsws = 0.037586
+ cjsws = {8.643094E-11*sw_func_nsd_pw_cj} cjswgs = {5.47776E-11*sw_func_nsd_pw_cj} mjswgs = 0.78692
+ pbs = 0.72468 pbsws = 0.29067 pbswgs = 0.54958
+ xrcrg1 = 12 xrcrg2 = 1 rbpb = 50
+ rbpd = 50 rbps = 50 rbdb = 50
+ rbsb = 50 gbmin = 1E-12 tnom = 30
+ ute = -1.068402 lute = -7.987541E-8 kt1 = -0.440127
+ lkt1 = 3.101958E-8 kt1l = 0 kt2 = -0.019151
+ ua1 = -1.43283E-9 lua1 = 1.539657E-15 ub1 = 1.705328E-18
+ lub1 = -1.409046E-24 wub1 = 7.250457E-23 pub1 = -3.240853E-29
+ uc1 = -5.9821E-11 at = -1.248544E5 lat = 6.87708E-2
+ wat = 1.643989 pat = -7.348402E-7 prt = 0
+ njs = 1.0773 xtis = 0.76 tpb = 1.344E-3
+ tpbsw = 9.9005E-4 tpbswg = 0 tcj = 6.7434E-4
+ tcjsw = 2.493E-4 tcjswg = 0 tvoff = 0
+ tvfbsdoff = 0 saref = 2.41E-6 sbref = 2.41E-6
+ wlod = 0 ku0 = -4.5E-8 kvsat = 0.3
+ kvth0 = 1.1E-8 tku0 = 0 llodku0 = 0
+ wlodku0 = 1 llodvth = 0 wlodvth = 1
+ lku0 = 0 wku0 = 2E-7 pku0 = 0
+ lkvth0 = 0 wkvth0 = 6.5E-7 pkvth0 = 0
+ stk2 = 0 lodk2 = 1 steta0 = 0
+ lodeta0 = 1

.model nhv_model.15 nmos
+ level = 54 lmin = 8E-6 lmax = 2.02E-5 wmin = 7E-6
+ wmax = 1.5E-5 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 1.16E-8
+ toxm = 1.16E-8 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 1E23 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {2.1346E-8+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {7.6507E-8-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = -4.1292E-9 dwb = -1.6944E-9 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = 0.78882 k1 = 0.88325
+ k2 = -0.039667 k3 = -0.884 k3b = 0.43
+ w0 = 0 lpe0 = 2.5E-8 lpeb = -2.182E-7
+ vbm = -3 dvtp0 = 0 dvtp1 = 0
+ dvt0 = 0 dvt1 = 0.53 dvt2 = -0.19251
+ dvt0w = 0.16 dvt1w = 6.9091E6 dvt2w = -0.036016
+ vfbsdoff = 0 u0 = 4.21082E-2 ua = -5.92431E-11
+ ub = 1.71671E-18 uc = 6.6204E-11 ud = 0
+ up = 0 lp = 1 eu = 1.67
+ vsat = 1.0566E5 a0 = 0.942599 ags = 0.149418
+ b0 = 3.2933E-8 b1 = 0 keta = -0.02132
+ a1 = 0 a2 = 0.659726 rdsw = 724.62
+ rdswmin = 0 rdw = 0 rdwmin = 0
+ rsw = 0 rswmin = 0 prwb = 0.05626
+ prwg = 0.048 wr = 1 voff = -0.20613
+ voffl = -4.257949E-7 minv = 0 nfactor = 0.96538
+ eta0 = 0.032 etab = -0.01932 dsub = 0.504
+ cit = -8E-4 cdsc = 0 cdscb = 0
+ cdscd = 0 pclm = 0.33405 pdiblc1 = 0.21098
+ pdiblc2 = 2E-4 pdiblcb = -0.26831 drout = 0.36075
+ pscbe1 = 9.3731E8 pscbe2 = 1.68E-6 pvag = 1.99
+ delta = 0.0246 fprout = 10.125 pdits = 0
+ pditsl = 0 pditsd = 0 lambda = 0
+ vtl = 0 lc = 5E-9 xn = 3
+ alpha0 = 1.4467E-5 alpha1 = 0 beta0 = 24
+ aigbacc = 1 bigbacc = 0 cigbacc = 0
+ nigbacc = 1 aigbinv = 0.35 bigbinv = 0.03
+ cigbinv = 6E-3 eigbinv = 1.1 nigbinv = 3
+ aigc = 0.43 bigc = 0.054 cigc = 0.075
+ aigsd = 0.43 bigsd = 0.054 cigsd = 0.075
+ dlcig = 0 nigc = 1 poxedge = 1
+ pigcd = 1 ntox = 1 toxref = 1.16E-8
+ agidl = 5.06E-11 bgidl = 1.058E9 cgidl = 4E3
+ egidl = 0.8 noia = 2.6E41 noib = 0
+ noic = 0 em = 4.1E7 af = 1
+ ef = 0.89 kf = 0 lintnoi = 0
+ tnoia = 7.5E6 tnoib = 7.2E6 ntnoi = 1
+ rnoia = 0.794 rnoib = 0.38 xpart = 0
+ cgso = {2.754679E-10/sw_func_tox_hv_ratio} cgdo = {2.754679E-10/sw_func_tox_hv_ratio} cgbo = {0/sw_func_tox_hv_ratio}
+ ckappas = 0.6 cf = 0 clc = 1E-7
+ cle = 0.6 dlc = 6.5995E-8 dwc = 0
+ vfbcv = -1 noff = 4 voffcv = -0.4104
+ acde = 0.4176 moin = 15 cgsl = {4.49025E-11/sw_func_tox_hv_ratio}
+ cgdl = {4.49025E-11/sw_func_tox_hv_ratio} ijthsrev = 0.1 ijthsfwd = 0.1
+ xjbvs = 1 bvs = 12.636 jss = 3.75E-4
+ jsws = 5.84E-11 cjs = {8.310E-04*sw_func_nsd_pw_cj} mjs = 0.295
+ mjsws = 0.037586 cjsws = {8.643094E-11*sw_func_nsd_pw_cj} cjswgs = {5.47776E-11*sw_func_nsd_pw_cj}
+ mjswgs = 0.78692 pbs = 0.72468 pbsws = 0.29067
+ pbswgs = 0.54958 xrcrg1 = 12 xrcrg2 = 1
+ rbpb = 50 rbpd = 50 rbps = 50
+ rbdb = 50 rbsb = 50 gbmin = 1E-12
+ tnom = 30 ute = -1.2986 kt1 = -0.40273
+ kt1l = 0 kt2 = -0.019151 ua1 = 3.0044E-9
+ ub1 = -3.7525E-18 uc1 = -5.9821E-11 at = 1.6E5
+ prt = 0 njs = 1.0773 xtis = 0.76
+ tpb = 1.344E-3 tpbsw = 9.9005E-4 tpbswg = 0
+ tcj = 6.7434E-4 tcjsw = 2.493E-4 tcjswg = 0
+ tvoff = 0 tvfbsdoff = 0 saref = 3E-6
+ sbref = 3E-6 wlod = 0 ku0 = -4.5E-8
+ kvsat = 0.3 kvth0 = 1.1E-8 tku0 = 0
+ llodku0 = 0 wlodku0 = 1 llodvth = 0
+ wlodvth = 1 lku0 = 0 wku0 = 2E-7
+ pku0 = 0 lkvth0 = 0 wkvth0 = 6.5E-7
+ pkvth0 = 0 stk2 = 0 lodk2 = 1
+ steta0 = 0 lodeta0 = 1

.model nhv_model.16 nmos
+ level = 54 lmin = 4E-6 lmax = 8E-6 wmin = 7E-6
+ wmax = 1.5E-5 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 1.16E-8
+ toxm = 1.16E-8 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 1E23 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {2.1346E-8+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {7.6507E-8-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = -4.1292E-9 dwb = -1.6944E-9 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = 0.783367 lvth0 = 4.279042E-8
+ k1 = 0.88325 k2 = -4.10016E-2 lk2 = 1.047271E-8
+ k3 = -0.884 k3b = 0.43 w0 = 0
+ lpe0 = 2.5E-8 lpeb = -2.182E-7 vbm = -3
+ dvtp0 = 0 dvtp1 = 0 dvt0 = 0
+ dvt1 = 0.53 dvt2 = -0.19251 dvt0w = 0.16
+ dvt1w = 6.9091E6 dvt2w = -0.036016 vfbsdoff = 0
+ u0 = 4.15573E-2 lu0 = 4.322814E-9 ua = -1.016037E-10
+ lua = 3.324031E-16 ub = 1.752362E-18 lub = -2.797603E-25
+ uc = 6.6204E-11 ud = 0 up = 0
+ lp = 1 eu = 1.67 vsat = 1.104687E5
+ lvsat = -3.77341E-2 a0 = 1.033611 la0 = -7.141721E-7
+ ags = 0.152066 lags = -2.078241E-8 b0 = 3.2933E-8
+ b1 = 0 keta = -1.72682E-2 lketa = -3.179472E-8
+ a1 = 0 a2 = 0.659726 rdsw = 724.62
+ rdswmin = 0 rdw = 0 rdwmin = 0
+ rsw = 0 rswmin = 0 prwb = 0.05626
+ prwg = 0.048 wr = 1 voff = -0.20613
+ voffl = -4.257949E-7 minv = 0 nfactor = 1.012092
+ lnfactor = -3.665486E-7 eta0 = 0.032 etab = -0.01932
+ dsub = 0.504 cit = -8E-4 cdsc = 0
+ cdscb = 0 cdscd = 0 pclm = 0.259909
+ lpclm = 5.817837E-7 pdiblc1 = 0.21098 pdiblc2 = 2E-4
+ pdiblcb = -0.26831 drout = 0.36075 pscbe1 = 9.3731E8
+ pscbe2 = 1.68E-6 pvag = 1.99 delta = 0.0246
+ fprout = 10.125 pdits = 0 pditsl = 0
+ pditsd = 0 lambda = 0 vtl = 0
+ lc = 5E-9 xn = 3 alpha0 = 1.4467E-5
+ alpha1 = 0 beta0 = 21.499459 lbeta0 = 1.962171E-5
+ aigbacc = 1 bigbacc = 0 cigbacc = 0
+ nigbacc = 1 aigbinv = 0.35 bigbinv = 0.03
+ cigbinv = 6E-3 eigbinv = 1.1 nigbinv = 3
+ aigc = 0.43 bigc = 0.054 cigc = 0.075
+ aigsd = 0.43 bigsd = 0.054 cigsd = 0.075
+ dlcig = 0 nigc = 1 poxedge = 1
+ pigcd = 1 ntox = 1 toxref = 1.16E-8
+ agidl = 5.06E-11 bgidl = 1.058E9 cgidl = 4E3
+ egidl = 0.8 noia = 2.6E41 noib = 0
+ noic = 0 em = 4.1E7 af = 1
+ ef = 0.89 kf = 0 lintnoi = 0
+ tnoia = 7.5E6 tnoib = 7.2E6 ntnoi = 1
+ rnoia = 0.794 rnoib = 0.38 xpart = 0
+ cgso = {2.754679E-10/sw_func_tox_hv_ratio} cgdo = {2.754679E-10/sw_func_tox_hv_ratio} cgbo = {0/sw_func_tox_hv_ratio}
+ ckappas = 0.6 cf = 0 clc = 1E-7
+ cle = 0.6 dlc = 6.5995E-8 dwc = 0
+ vfbcv = -1 noff = 4 voffcv = -0.4104
+ acde = 0.4176 moin = 15 cgsl = {4.49025E-11/sw_func_tox_hv_ratio}
+ cgdl = {4.49025E-11/sw_func_tox_hv_ratio} ijthsrev = 0.1 ijthsfwd = 0.1
+ xjbvs = 1 bvs = 12.636 jss = 3.75E-4
+ jsws = 5.84E-11 cjs = {8.310E-04*sw_func_nsd_pw_cj} mjs = 0.295
+ mjsws = 0.037586 cjsws = {8.643094E-11*sw_func_nsd_pw_cj} cjswgs = {5.47776E-11*sw_func_nsd_pw_cj}
+ mjswgs = 0.78692 pbs = 0.72468 pbsws = 0.29067
+ pbswgs = 0.54958 xrcrg1 = 12 xrcrg2 = 1
+ rbpb = 50 rbpd = 50 rbps = 50
+ rbdb = 50 rbsb = 50 gbmin = 1E-12
+ tnom = 30 ute = -1.33707 lute = 3.018725E-7
+ kt1 = -0.414271 lkt1 = 9.056174E-8 kt1l = 0
+ kt2 = -0.019151 ua1 = 3.0044E-9 ub1 = -3.7525E-18
+ uc1 = -5.9821E-11 at = 2.369397E5 lat = -0.603745
+ prt = 0 njs = 1.0773 xtis = 0.76
+ tpb = 1.344E-3 tpbsw = 9.9005E-4 tpbswg = 0
+ tcj = 6.7434E-4 tcjsw = 2.493E-4 tcjswg = 0
+ tvoff = 0 tvfbsdoff = 0 saref = 3E-6
+ sbref = 3E-6 wlod = 0 ku0 = -4.5E-8
+ kvsat = 0.3 kvth0 = 1.1E-8 tku0 = 0
+ llodku0 = 0 wlodku0 = 1 llodvth = 0
+ wlodvth = 1 lku0 = 0 wku0 = 2E-7
+ pku0 = 0 lkvth0 = 0 wkvth0 = 6.5E-7
+ pkvth0 = 0 stk2 = 0 lodk2 = 1
+ steta0 = 0 lodeta0 = 1

.model nhv_model.17 nmos
+ level = 54 lmin = 2E-6 lmax = 4E-6 wmin = 7E-6
+ wmax = 1.5E-5 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 1.16E-8
+ toxm = 1.16E-8 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 1E23 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {2.1346E-8+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {7.6507E-8-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = -4.1292E-9 dwb = -1.6944E-9 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = 0.799231 lvth0 = -1.823938E-8
+ k1 = 0.88325 k2 = -4.25688E-2 lk2 = 1.650177E-8
+ k3 = -0.884 k3b = 0.43 w0 = 0
+ lpe0 = 2.5E-8 lpeb = -2.182E-7 vbm = -3
+ dvtp0 = 0 dvtp1 = 0 dvt0 = 0
+ dvt1 = 0.53 dvt2 = -0.19251 dvt0w = 0.16
+ dvt1w = 6.9091E6 dvt2w = -0.036016 vfbsdoff = 0
+ u0 = 4.27638E-2 lu0 = -3.18674E-10 ua = 1.059937E-10
+ lua = -4.662212E-16 ub = 1.549686E-18 lub = 4.99931E-25
+ uc = 6.6204E-11 ud = 0 up = 0
+ lp = 1 eu = 1.67 vsat = 9.377998E4
+ lvsat = 2.64674E-2 a0 = 0.476534 la0 = 1.428898E-6
+ ags = 0.119435 lags = 1.047503E-7 b0 = 3.2933E-8
+ b1 = 0 keta = -3.92681E-2 lketa = 5.283878E-8
+ a1 = 0 a2 = 0.659726 rdsw = 724.62
+ rdswmin = 0 rdw = 0 rdwmin = 0
+ rsw = 0 rswmin = 0 prwb = 0.05626
+ prwg = 0.048 wr = 1 voff = -0.20613
+ voffl = -4.257949E-7 minv = 0 nfactor = 0.961332
+ lnfactor = -1.71274E-7 eta0 = 0.032 etab = -0.01932
+ dsub = 0.504 cit = -8E-4 cdsc = 0
+ cdscb = 0 cdscd = 0 pclm = 0.600982
+ lpclm = -7.303213E-7 pdiblc1 = 0.21098 pdiblc2 = 2E-4
+ pdiblcb = -0.26831 drout = 0.36075 pscbe1 = 9.3731E8
+ pscbe2 = 1.68E-6 pvag = 1.99 delta = 0.0246
+ fprout = 10.125 pdits = 0 pditsl = 0
+ pditsd = 0 lambda = 0 vtl = 0
+ lc = 5E-9 xn = 3 alpha0 = 1.4467E-5
+ alpha1 = 0 beta0 = 23.859073 lbeta0 = 1.054431E-5
+ aigbacc = 1 bigbacc = 0 cigbacc = 0
+ nigbacc = 1 aigbinv = 0.35 bigbinv = 0.03
+ cigbinv = 6E-3 eigbinv = 1.1 nigbinv = 3
+ aigc = 0.43 bigc = 0.054 cigc = 0.075
+ aigsd = 0.43 bigsd = 0.054 cigsd = 0.075
+ dlcig = 0 nigc = 1 poxedge = 1
+ pigcd = 1 ntox = 1 toxref = 1.16E-8
+ agidl = 5.06E-11 bgidl = 1.058E9 cgidl = 4E3
+ egidl = 0.8 noia = 2.6E41 noib = 0
+ noic = 0 em = 4.1E7 af = 1
+ ef = 0.89 kf = 0 lintnoi = 0
+ tnoia = 7.5E6 tnoib = 7.2E6 ntnoi = 1
+ rnoia = 0.794 rnoib = 0.38 xpart = 0
+ cgso = {2.754679E-10/sw_func_tox_hv_ratio} cgdo = {2.754679E-10/sw_func_tox_hv_ratio} cgbo = {0/sw_func_tox_hv_ratio}
+ ckappas = 0.6 cf = 0 clc = 1E-7
+ cle = 0.6 dlc = 6.5995E-8 dwc = 0
+ vfbcv = -1 noff = 4 voffcv = -0.4104
+ acde = 0.4176 moin = 15 cgsl = {4.49025E-11/sw_func_tox_hv_ratio}
+ cgdl = {4.49025E-11/sw_func_tox_hv_ratio} ijthsrev = 0.1 ijthsfwd = 0.1
+ xjbvs = 1 bvs = 12.636 jss = 3.75E-4
+ jsws = 5.84E-11 cjs = {8.310E-04*sw_func_nsd_pw_cj} mjs = 0.295
+ mjsws = 0.037586 cjsws = {8.643094E-11*sw_func_nsd_pw_cj} cjswgs = {5.47776E-11*sw_func_nsd_pw_cj}
+ mjswgs = 0.78692 pbs = 0.72468 pbsws = 0.29067
+ pbswgs = 0.54958 xrcrg1 = 12 xrcrg2 = 1
+ rbpb = 50 rbpd = 50 rbps = 50
+ rbdb = 50 rbsb = 50 gbmin = 1E-12
+ tnom = 30 ute = -1.22166 lute = -1.421066E-7
+ kt1 = -0.407353 lkt1 = 6.394796E-8 kt1l = 0
+ kt2 = -0.019151 ua1 = 3.0044E-9 ub1 = -3.7525E-18
+ uc1 = -5.9821E-11 at = 1.391036E5 lat = -0.227371
+ prt = 0 njs = 1.0773 xtis = 0.76
+ tpb = 1.344E-3 tpbsw = 9.9005E-4 tpbswg = 0
+ tcj = 6.7434E-4 tcjsw = 2.493E-4 tcjswg = 0
+ tvoff = 0 tvfbsdoff = 0 saref = 3E-6
+ sbref = 3E-6 wlod = 0 ku0 = -4.5E-8
+ kvsat = 0.3 kvth0 = 1.1E-8 tku0 = 0
+ llodku0 = 0 wlodku0 = 1 llodvth = 0
+ wlodvth = 1 lku0 = 0 wku0 = 2E-7
+ pku0 = 0 lkvth0 = 0 wkvth0 = 6.5E-7
+ pkvth0 = 0 stk2 = 0 lodk2 = 1
+ steta0 = 0 lodeta0 = 1

.model nhv_model.18 nmos
+ level = 54 lmin = 1E-6 lmax = 2E-6 wmin = 7E-6
+ wmax = 1.5E-5 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 1.16E-8
+ toxm = 1.16E-8 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 1E23 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {2.1346E-8+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {7.6507E-8-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = -4.1292E-9 dwb = -1.6944E-9 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = 0.774727 lvth0 = 2.701999E-8
+ wvth0 = 5.087856E-8 pvth0 = -9.397199E-14 k1 = 0.88325
+ k2 = -4.01544E-2 lk2 = 1.204241E-8 wk2 = -1.134577E-8
+ pk2 = 2.095547E-14 k3 = -0.884 k3b = 0.43
+ w0 = 0 lpe0 = 2.5E-8 lpeb = -2.182E-7
+ vbm = -3 dvtp0 = 0 dvtp1 = 0
+ dvt0 = 0 dvt1 = 0.53 dvt2 = -0.19251
+ dvt0w = 0.16 dvt1w = 6.9091E6 dvt2w = -0.036016
+ vfbsdoff = 0 u0 = 4.11832E-2 lu0 = 2.600652E-9
+ wu0 = 2.887011E-9 pu0 = -5.33227E-15 ua = -1.362862E-10
+ lua = -1.873361E-17 wua = -5.730614E-17 pua = 1.058436E-22
+ ub = 1.776248E-18 lub = 8.147357E-26 wub = 3.236925E-25
+ pub = -5.978556E-31 uc = 6.6204E-11 ud = 0
+ up = 0 lp = 1 eu = 1.67
+ vsat = 1.204553E5 lvsat = -2.28016E-2 wvsat = -4.65267E-2
+ pvsat = 8.593411E-8 a0 = 2.061458 la0 = -1.498436E-6
+ wa0 = -5.65247E-6 pa0 = 1.044003E-11 ags = 0.196716
+ lags = -3.798611E-8 wags = -8.193344E-8 pags = 1.513299E-13
+ b0 = 3.2933E-8 b1 = 0 keta = 1.54817E-2
+ lketa = -4.828339E-8 wketa = -1.81876E-7 pketa = 3.359224E-13
+ a1 = 0 a2 = 0.659726 rdsw = 724.62
+ rdswmin = 0 rdw = 0 rdwmin = 0
+ rsw = 0 rswmin = 0 prwb = 0.05626
+ prwg = 0.048 wr = 1 voff = -0.20613
+ voffl = -4.257949E-7 minv = 0 nfactor = 0.899606
+ lnfactor = -5.72678E-8 wnfactor = 3.10692E-8 pnfactor = -5.738437E-14
+ eta0 = 0.032 etab = -0.01932 dsub = 0.504
+ cit = -8E-4 cdsc = 0 cdscb = 0
+ cdscd = 0 pclm = 0.380662 lpclm = -3.233917E-7
+ wpclm = -4.246564E-6 ppclm = 7.843345E-12 pdiblc1 = 0.21098
+ pdiblc2 = 2E-4 pdiblcb = -0.26831 drout = 0.36075
+ pscbe1 = 9.3731E8 pscbe2 = 1.68E-6 pvag = 1.99
+ delta = 0.0246 fprout = 10.125 pdits = 0
+ pditsl = 0 pditsd = 0 lambda = 0
+ vtl = 0 lc = 5E-9 xn = 3
+ alpha0 = 1.361476E-5 lalpha0 = 1.574071E-12 walpha0 = 1.274718E-11
+ palpha0 = -2.354387E-17 alpha1 = 0 beta0 = 27.266025
+ lbeta0 = 4.251715E-6 wbeta0 = -3.029798E-6 pbeta0 = 5.595994E-12
+ aigbacc = 1 bigbacc = 0 cigbacc = 0
+ nigbacc = 1 aigbinv = 0.35 bigbinv = 0.03
+ cigbinv = 6E-3 eigbinv = 1.1 nigbinv = 3
+ aigc = 0.43 bigc = 0.054 cigc = 0.075
+ aigsd = 0.43 bigsd = 0.054 cigsd = 0.075
+ dlcig = 0 nigc = 1 poxedge = 1
+ pigcd = 1 ntox = 1 toxref = 1.16E-8
+ agidl = 5.06E-11 bgidl = 1.058E9 cgidl = 4E3
+ egidl = 0.8 noia = 2.6E41 noib = 0
+ noic = 0 em = 4.1E7 af = 1
+ ef = 0.89 kf = 0 lintnoi = 0
+ tnoia = 7.5E6 tnoib = 7.2E6 ntnoi = 1
+ rnoia = 0.794 rnoib = 0.38 xpart = 0
+ cgso = {2.754679E-10/sw_func_tox_hv_ratio} cgdo = {2.754679E-10/sw_func_tox_hv_ratio} cgbo = {0/sw_func_tox_hv_ratio}
+ ckappas = 0.6 cf = 0 clc = 1E-7
+ cle = 0.6 dlc = 6.5995E-8 dwc = 0
+ vfbcv = -1 noff = 4 voffcv = -0.4104
+ acde = 0.4176 moin = 15 cgsl = {4.49025E-11/sw_func_tox_hv_ratio}
+ cgdl = {4.49025E-11/sw_func_tox_hv_ratio} ijthsrev = 0.1 ijthsfwd = 0.1
+ xjbvs = 1 bvs = 12.636 jss = 3.75E-4
+ jsws = 5.84E-11 cjs = {8.310E-04*sw_func_nsd_pw_cj} mjs = 0.295
+ mjsws = 0.037586 cjsws = {8.643094E-11*sw_func_nsd_pw_cj} cjswgs = {5.47776E-11*sw_func_nsd_pw_cj}
+ mjswgs = 0.78692 pbs = 0.72468 pbsws = 0.29067
+ pbswgs = 0.54958 xrcrg1 = 12 xrcrg2 = 1
+ rbpb = 50 rbpd = 50 rbps = 50
+ rbdb = 50 rbsb = 50 gbmin = 1E-12
+ tnom = 30 ute = -1.2986 kt1 = -0.388566
+ lkt1 = 2.924848E-8 wkt1 = 1.101745E-7 pkt1 = -2.034907E-13
+ kt1l = 0 kt2 = -0.019151 ua1 = 3.0044E-9
+ ub1 = -4.22789E-18 lub1 = 8.780393E-25 wub1 = 3.307437E-24
+ pub1 = -6.10879E-30 uc1 = -5.9821E-11 at = 9.224112E3
+ lat = 0.012515 prt = 0 njs = 1.0773
+ xtis = 0.76 tpb = 1.344E-3 tpbsw = 9.9005E-4
+ tpbswg = 0 tcj = 6.7434E-4 tcjsw = 2.493E-4
+ tcjswg = 0 tvoff = 0 tvfbsdoff = 0
+ saref = 3E-6 sbref = 3E-6 wlod = 0
+ ku0 = -4.5E-8 kvsat = 0.3 kvth0 = 1.1E-8
+ tku0 = 0 llodku0 = 0 wlodku0 = 1
+ llodvth = 0 wlodvth = 1 lku0 = 0
+ wku0 = 2E-7 pku0 = 0 lkvth0 = 0
+ wkvth0 = 6.5E-7 pkvth0 = 0 stk2 = 0
+ lodk2 = 1 steta0 = 0 lodeta0 = 1

.model nhv_model.19 nmos
+ level = 54 lmin = 8E-7 lmax = 1E-6 wmin = 7E-6
+ wmax = 1.5E-5 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 1.16E-8
+ toxm = 1.16E-8 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 1E23 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {2.1346E-8+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {7.6507E-8-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = -4.1292E-9 dwb = -1.6944E-9 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = 0.807288 lvth0 = -5.592384E-10
+ wvth0 = -2.543928E-7 pvth0 = 1.645886E-13 k1 = 0.88325
+ k2 = -3.88774E-2 lk2 = 1.09608E-8 wk2 = 5.672883E-8
+ pk2 = -3.670276E-14 k3 = -0.884 k3b = 0.43
+ w0 = 0 lpe0 = 2.5E-8 lpeb = -2.182E-7
+ vbm = -3 dvtp0 = 0 dvtp1 = 0
+ dvt0 = 0 dvt1 = 0.53 dvt2 = -0.19251
+ dvt0w = 0.16 dvt1w = 6.9091E6 dvt2w = -0.036016
+ vfbsdoff = 0 u0 = 4.55329E-2 lu0 = -1.083445E-9
+ wu0 = -1.443506E-8 pu0 = 9.33928E-15 ua = -1.913677E-10
+ lua = 2.791963E-17 wua = 2.865307E-16 pua = -1.853814E-22
+ ub = 1.536528E-18 lub = 2.845135E-25 wub = -1.618463E-24
+ pub = 1.047123E-30 uc = 6.6204E-11 ud = 0
+ up = 0 lp = 1 eu = 1.67
+ vsat = 8.227786E4 lvsat = 9.53414E-3 wvsat = 0.232633
+ pvsat = -1.505105E-7 a0 = -2.392288 la0 = 2.273825E-6
+ wa0 = 2.826235E-5 pa0 = -1.828534E-11 ags = 0.124748
+ lags = 2.296899E-8 wags = 4.096672E-7 pags = -2.650489E-13
+ b0 = 3.2933E-8 b1 = 0 keta = -0.141369
+ lketa = 8.456663E-8 wketa = 9.0938E-7 pketa = -5.883561E-13
+ a1 = 0 a2 = 0.659726 rdsw = 724.62
+ rdswmin = 0 rdw = 0 rdwmin = 0
+ rsw = 0 rswmin = 0 prwb = 0.05626
+ prwg = 0.048 wr = 1 voff = -0.20613
+ voffl = -4.257949E-7 minv = 0 nfactor = 0.864835
+ lnfactor = -2.781711E-8 wnfactor = -1.55346E-7 pnfactor = 1.005067E-13
+ eta0 = 0.032 etab = -0.01932 dsub = 0.504
+ cit = -8E-4 cdsc = 0 cdscb = 0
+ cdscd = 0 pclm = -3.329744 lpclm = 2.81927E-6
+ wpclm = 2.123282E-5 ppclm = -1.373734E-11 pdiblc1 = 0.21098
+ pdiblc2 = 2E-4 pdiblcb = -0.26831 drout = 0.36075
+ pscbe1 = 9.3731E8 pscbe2 = 1.68E-6 pvag = 1.99
+ delta = 0.0246 fprout = 10.125 pdits = 0
+ pditsl = 0 pditsd = 0 lambda = 0
+ vtl = 0 lc = 5E-9 xn = 3
+ alpha0 = 9.369537E-6 lalpha0 = 5.169718E-12 walpha0 = -6.373592E-11
+ palpha0 = 4.123625E-17 alpha1 = 0 beta0 = 21.946497
+ lbeta0 = 8.757281E-6 wbeta0 = 1.514899E-5 pbeta0 = -9.801183E-12
+ aigbacc = 1 bigbacc = 0 cigbacc = 0
+ nigbacc = 1 aigbinv = 0.35 bigbinv = 0.03
+ cigbinv = 6E-3 eigbinv = 1.1 nigbinv = 3
+ aigc = 0.43 bigc = 0.054 cigc = 0.075
+ aigsd = 0.43 bigsd = 0.054 cigsd = 0.075
+ dlcig = 0 nigc = 1 poxedge = 1
+ pigcd = 1 ntox = 1 toxref = 1.16E-8
+ agidl = 5.06E-11 bgidl = 1.058E9 cgidl = 4E3
+ egidl = 0.8 noia = 2.6E41 noib = 0
+ noic = 0 em = 4.1E7 af = 1
+ ef = 0.89 kf = 0 lintnoi = 0
+ tnoia = 7.5E6 tnoib = 7.2E6 ntnoi = 1
+ rnoia = 0.794 rnoib = 0.38 xpart = 0
+ cgso = {2.754679E-10/sw_func_tox_hv_ratio} cgdo = {2.754679E-10/sw_func_tox_hv_ratio} cgbo = {0/sw_func_tox_hv_ratio}
+ ckappas = 0.6 cf = 0 clc = 1E-7
+ cle = 0.6 dlc = 6.5995E-8 dwc = 0
+ vfbcv = -1 noff = 4 voffcv = -0.4104
+ acde = 0.4176 moin = 15 cgsl = {4.49025E-11/sw_func_tox_hv_ratio}
+ cgdl = {4.49025E-11/sw_func_tox_hv_ratio} ijthsrev = 0.1 ijthsfwd = 0.1
+ xjbvs = 1 bvs = 12.636 jss = 3.75E-4
+ jsws = 5.84E-11 cjs = {8.310E-04*sw_func_nsd_pw_cj} mjs = 0.295
+ mjsws = 0.037586 cjsws = {8.643094E-11*sw_func_nsd_pw_cj} cjswgs = {5.47776E-11*sw_func_nsd_pw_cj}
+ mjswgs = 0.78692 pbs = 0.72468 pbsws = 0.29067
+ pbswgs = 0.54958 xrcrg1 = 12 xrcrg2 = 1
+ rbpb = 50 rbpd = 50 rbps = 50
+ rbdb = 50 rbsb = 50 gbmin = 1E-12
+ tnom = 30 ute = -1.465199 lute = 1.411069E-7
+ kt1 = -0.300021 lkt1 = -4.574779E-8 wkt1 = -5.508723E-7
+ pkt1 = 3.564067E-13 kt1l = 0 kt2 = -0.019151
+ ua1 = 6.215715E-9 lua1 = -2.719939E-15 ub1 = -8.833679E-18
+ lub1 = 4.779078E-24 wub1 = -1.653719E-23 pub1 = 1.069933E-29
+ uc1 = -5.9821E-11 at = 7.82535E3 lat = 1.36997E-2
+ prt = 0 njs = 1.0773 xtis = 0.76
+ tpb = 1.344E-3 tpbsw = 9.9005E-4 tpbswg = 0
+ tcj = 6.7434E-4 tcjsw = 2.493E-4 tcjswg = 0
+ tvoff = 0 tvfbsdoff = 0 saref = 2.81E-6
+ sbref = 2.81E-6 wlod = 0 ku0 = -4.5E-8
+ kvsat = 0.3 kvth0 = 1.1E-8 tku0 = 0
+ llodku0 = 0 wlodku0 = 1 llodvth = 0
+ wlodvth = 1 lku0 = 0 wku0 = 2E-7
+ pku0 = 0 lkvth0 = 0 wkvth0 = 6.5E-7
+ pkvth0 = 0 stk2 = 0 lodk2 = 1
+ steta0 = 0 lodeta0 = 1

.model nhv_model.20 nmos
+ level = 54 lmin = 6E-7 lmax = 8E-7 wmin = 7E-6
+ wmax = 1.5E-5 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 1.16E-8
+ toxm = 1.16E-8 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 1E23 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {2.1346E-8+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {7.6507E-8-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = -4.1292E-9 dwb = -1.6944E-9 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = 0.806424 k1 = 0.88325
+ k2 = -2.19361E-2 k3 = -0.884 k3b = 0.43
+ w0 = 0 lpe0 = 2.5E-8 lpeb = -2.182E-7
+ vbm = -3 dvtp0 = 0 dvtp1 = 0
+ dvt0 = 0 dvt1 = 0.53 dvt2 = -0.19251
+ dvt0w = 0.16 dvt1w = 6.9091E6 dvt2w = -0.036016
+ vfbsdoff = 0 u0 = 4.38583E-2 ua = -1.482143E-10
+ ub = 1.97628E-18 uc = 6.6204E-11 ud = 0
+ up = 0 lp = 1 eu = 1.67
+ vsat = 9.70141E4 a0 = 1.1222 ags = 0.16025
+ b0 = 3.2933E-8 b1 = 0 keta = -0.01066
+ a1 = 0 a2 = 0.659726 rdsw = 724.62
+ rdswmin = 0 rdw = 0 rdwmin = 0
+ rsw = 0 rswmin = 0 prwb = 0.05626
+ prwg = 0.048 wr = 1 voff = -0.20613
+ voffl = -4.257949E-7 minv = 0 nfactor = 0.82184
+ eta0 = 0.032 etab = -0.01932 dsub = 0.504
+ cit = -8E-4 cdsc = 0 cdscb = 0
+ cdscd = 0 pclm = 1.0278 pdiblc1 = 0.21098
+ pdiblc2 = 2E-4 pdiblcb = -0.26831 drout = 0.36075
+ pscbe1 = 9.3731E8 pscbe2 = 1.68E-6 pvag = 1.99
+ delta = 0.0246 fprout = 10.125 pdits = 0
+ pditsl = 0 pditsd = 0 lambda = 0
+ vtl = 0 lc = 5E-9 xn = 3
+ alpha0 = 1.736E-5 alpha1 = 0 beta0 = 35.482
+ aigbacc = 1 bigbacc = 0 cigbacc = 0
+ nigbacc = 1 aigbinv = 0.35 bigbinv = 0.03
+ cigbinv = 6E-3 eigbinv = 1.1 nigbinv = 3
+ aigc = 0.43 bigc = 0.054 cigc = 0.075
+ aigsd = 0.43 bigsd = 0.054 cigsd = 0.075
+ dlcig = 0 nigc = 1 poxedge = 1
+ pigcd = 1 ntox = 1 toxref = 1.16E-8
+ agidl = 5.06E-11 bgidl = 1.058E9 cgidl = 4E3
+ egidl = 0.8 noia = 2.6E41 noib = 0
+ noic = 0 em = 4.1E7 af = 1
+ ef = 0.89 kf = 0 lintnoi = 0
+ tnoia = 7.5E6 tnoib = 7.2E6 ntnoi = 1
+ rnoia = 0.794 rnoib = 0.38 xpart = 0
+ cgso = {2.754679E-10/sw_func_tox_hv_ratio} cgdo = {2.754679E-10/sw_func_tox_hv_ratio} cgbo = {0/sw_func_tox_hv_ratio}
+ ckappas = 0.6 cf = 0 clc = 1E-7
+ cle = 0.6 dlc = 6.5995E-8 dwc = 0
+ vfbcv = -1 noff = 4 voffcv = -0.4104
+ acde = 0.4176 moin = 15 cgsl = {4.49025E-11/sw_func_tox_hv_ratio}
+ cgdl = {4.49025E-11/sw_func_tox_hv_ratio} ijthsrev = 0.1 ijthsfwd = 0.1
+ xjbvs = 1 bvs = 12.636 jss = 3.75E-4
+ jsws = 5.84E-11 cjs = {8.310E-04*sw_func_nsd_pw_cj} mjs = 0.295
+ mjsws = 0.037586 cjsws = {8.643094E-11*sw_func_nsd_pw_cj} cjswgs = {5.47776E-11*sw_func_nsd_pw_cj}
+ mjswgs = 0.78692 pbs = 0.72468 pbsws = 0.29067
+ pbswgs = 0.54958 xrcrg1 = 12 xrcrg2 = 1
+ rbpb = 50 rbpd = 50 rbps = 50
+ rbdb = 50 rbsb = 50 gbmin = 1E-12
+ tnom = 30 ute = -1.2471 kt1 = -0.37073
+ kt1l = 0 kt2 = -0.019151 ua1 = 2.0117E-9
+ ub1 = -1.447E-18 uc1 = -5.9821E-11 at = 2.9E4
+ prt = 0 njs = 1.0773 xtis = 0.76
+ tpb = 1.344E-3 tpbsw = 9.9005E-4 tpbswg = 0
+ tcj = 6.7434E-4 tcjsw = 2.493E-4 tcjswg = 0
+ tvoff = 0 tvfbsdoff = 0 saref = 2.41E-6
+ sbref = 2.41E-6 wlod = 0 ku0 = -4.5E-8
+ kvsat = 0.3 kvth0 = 1.1E-8 tku0 = 0
+ llodku0 = 0 wlodku0 = 1 llodvth = 0
+ wlodvth = 1 lku0 = 0 wku0 = 2E-7
+ pku0 = 0 lkvth0 = 0 wkvth0 = 6.5E-7
+ pkvth0 = 0 stk2 = 0 lodk2 = 1
+ steta0 = 0 lodeta0 = 1

.model nhv_model.21 nmos
+ level = 54 lmin = 5E-7 lmax = 6E-7 wmin = 7E-6
+ wmax = 1.5E-5 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 1.16E-8
+ toxm = 1.16E-8 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 1E23 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {2.1346E-8+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {7.6507E-8-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = -4.1292E-9 dwb = -1.6944E-9 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = 0.758815 lvth0 = 2.128049E-8
+ wvth0 = 4.731537E-7 pvth0 = -2.114931E-13 k1 = 0.88325
+ k2 = 2.13933E-2 lk2 = -1.936763E-8 wk2 = -3.235752E-8
+ pk2 = 1.446336E-14 k3 = -0.884 k3b = 0.43
+ w0 = 0 lpe0 = 2.5E-8 lpeb = -2.182E-7
+ vbm = -3 dvtp0 = 0 dvtp1 = 0
+ dvt0 = 0 dvt1 = 0.53 dvt2 = -0.19251
+ dvt0w = 0.16 dvt1w = 6.9091E6 dvt2w = -0.036016
+ vfbsdoff = 0 u0 = 2.12034E-2 lu0 = 1.012644E-8
+ wu0 = 3.263284E-8 pu0 = -1.458642E-14 ua = -1.220513E-10
+ lua = -1.169448E-17 wua = -1.332404E-16 pua = 5.955659E-23
+ ub = -2.169597E-18 lub = 1.853149E-24 wub = 5.092168E-24
+ pub = -2.276128E-30 uc = 6.6204E-11 ud = 0
+ up = 0 lp = 1 eu = 1.67
+ vsat = 6.617771E4 lvsat = 1.37834E-2 wvsat = 2.49698E-2
+ pvsat = -1.116114E-8 a0 = 1.1222 ags = 0.16025
+ b0 = 3.2933E-8 b1 = 0 keta = -0.01066
+ a1 = 0 a2 = 0.659726 rdsw = 724.62
+ rdswmin = 0 rdw = 0 rdwmin = 0
+ rsw = 0 rswmin = 0 prwb = 0.05626
+ prwg = 0.048 wr = 1 voff = -0.20613
+ voffl = -4.257949E-7 minv = 0 nfactor = 1.19894
+ lnfactor = -1.685584E-7 wnfactor = -1.396036E-6 pnfactor = 6.240085E-13
+ eta0 = 0.032 etab = -0.01932 dsub = 0.504
+ cit = -8E-4 cdsc = 0 cdscb = 0
+ cdscd = 0 pclm = 1.46987 lpclm = -1.975991E-7
+ wpclm = -9.279824E-6 ppclm = 4.147951E-12 pdiblc1 = 0.21098
+ pdiblc2 = 2E-4 pdiblcb = -0.26831 drout = 0.36075
+ pscbe1 = 9.3731E8 pscbe2 = 1.68E-6 pvag = 1.99
+ delta = 0.0246 fprout = 10.125 pdits = 0
+ pditsl = 0 pditsd = 0 lambda = 0
+ vtl = 0 lc = 5E-9 xn = 3
+ alpha0 = 2.73983E-5 lalpha0 = -4.486982E-12 alpha1 = 0
+ beta0 = 30.353547 lbeta0 = 2.292347E-6 aigbacc = 1
+ bigbacc = 0 cigbacc = 0 nigbacc = 1
+ aigbinv = 0.35 bigbinv = 0.03 cigbinv = 6E-3
+ eigbinv = 1.1 nigbinv = 3 aigc = 0.43
+ bigc = 0.054 cigc = 0.075 aigsd = 0.43
+ bigsd = 0.054 cigsd = 0.075 dlcig = 0
+ nigc = 1 poxedge = 1 pigcd = 1
+ ntox = 1 toxref = 1.16E-8 agidl = 5.06E-11
+ bgidl = 1.058E9 cgidl = 4E3 egidl = 0.8
+ noia = 2.6E41 noib = 0 noic = 0
+ em = 4.1E7 af = 1 ef = 0.89
+ kf = 0 lintnoi = 0 tnoia = 7.5E6
+ tnoib = 7.2E6 ntnoi = 1 rnoia = 0.794
+ rnoib = 0.38 xpart = 0 cgso = {2.754679E-10/sw_func_tox_hv_ratio}
+ cgdo = {2.754679E-10/sw_func_tox_hv_ratio} cgbo = {0/sw_func_tox_hv_ratio} ckappas = 0.6
+ cf = 0 clc = 1E-7 cle = 0.6
+ dlc = 6.5995E-8 dwc = 0 vfbcv = -1
+ noff = 4 voffcv = -0.4104 acde = 0.4176
+ moin = 15 cgsl = {4.49025E-11/sw_func_tox_hv_ratio} cgdl = {4.49025E-11/sw_func_tox_hv_ratio}
+ ijthsrev = 0.1 ijthsfwd = 0.1 xjbvs = 1
+ bvs = 12.636 jss = 3.75E-4 jsws = 5.84E-11
+ cjs = {8.310E-04*sw_func_nsd_pw_cj} mjs = 0.295 mjsws = 0.037586
+ cjsws = {8.643094E-11*sw_func_nsd_pw_cj} cjswgs = {5.47776E-11*sw_func_nsd_pw_cj} mjswgs = 0.78692
+ pbs = 0.72468 pbsws = 0.29067 pbswgs = 0.54958
+ xrcrg1 = 12 xrcrg2 = 1 rbpb = 50
+ rbpd = 50 rbps = 50 rbdb = 50
+ rbsb = 50 gbmin = 1E-12 tnom = 30
+ ute = -1.068402 lute = -7.987541E-8 kt1 = -0.440127
+ lkt1 = 3.101958E-8 kt1l = 0 kt2 = -0.019151
+ ua1 = -1.43283E-9 lua1 = 1.539657E-15 ub1 = 7.156284E-18
+ lub1 = -3.845548E-24 wub1 = -9.027066E-24 pub1 = 4.034972E-30
+ uc1 = -5.9821E-11 at = -1.996361E4 lat = 0.021886
+ wat = 7.51052E-2 pat = -3.357097E-8 prt = 0
+ njs = 1.0773 xtis = 0.76 tpb = 1.344E-3
+ tpbsw = 9.9005E-4 tpbswg = 0 tcj = 6.7434E-4
+ tcjsw = 2.493E-4 tcjswg = 0 tvoff = 0
+ tvfbsdoff = 0 saref = 2.41E-6 sbref = 2.41E-6
+ wlod = 0 ku0 = -4.5E-8 kvsat = 0.3
+ kvth0 = 1.1E-8 tku0 = 0 llodku0 = 0
+ wlodku0 = 1 llodvth = 0 wlodvth = 1
+ lku0 = 0 wku0 = 2E-7 pku0 = 0
+ lkvth0 = 0 wkvth0 = 6.5E-7 pkvth0 = 0
+ stk2 = 0 lodk2 = 1 steta0 = 0
+ lodeta0 = 1

.model nhv_model.22 nmos
+ level = 54 lmin = 8E-6 lmax = 2.02E-5 wmin = 5E-6
+ wmax = 7E-6 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 1.16E-8
+ toxm = 1.16E-8 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 1E23 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {2.1346E-8+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {7.6507E-8-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = -4.1292E-9 dwb = -1.6944E-9 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = 0.773931 wvth0 = 1.035893E-7
+ k1 = 0.88325 k2 = -3.90052E-2 wk2 = -4.604351E-9
+ k3 = -0.884 k3b = 0.43 w0 = 0
+ lpe0 = 2.5E-8 lpeb = -2.182E-7 vbm = -3
+ dvtp0 = 0 dvtp1 = 0 dvt0 = 0
+ dvt1 = 0.53 dvt2 = -0.19251 dvt0w = 0.16
+ dvt1w = 6.9091E6 dvt2w = -0.036016 vfbsdoff = 0
+ u0 = 4.12945E-2 wu0 = 5.661454E-9 ua = -3.776292E-10
+ wua = 2.21511E-15 ub = 2.154217E-18 wub = -3.043872E-24
+ uc = 6.6204E-11 ud = 0 up = 0
+ lp = 1 eu = 1.67 vsat = 1.192182E5
+ wvsat = -9.43288E-2 a0 = 1.229923 wa0 = -1.999E-6
+ ags = 0.169888 wags = -1.424176E-7 b0 = 3.2933E-8
+ b1 = 0 keta = -1.70294E-2 wketa = -2.985068E-8
+ a1 = 0 a2 = 0.659726 rdsw = 724.62
+ rdswmin = 0 rdw = 0 rdwmin = 0
+ rsw = 0 rswmin = 0 prwb = 0.05626
+ prwg = 0.048 wr = 1 voff = -0.20613
+ voffl = -4.257949E-7 minv = 0 nfactor = 0.908916
+ wnfactor = 3.928356E-7 eta0 = 0.032 etab = -0.01932
+ dsub = 0.504 cit = -8E-4 cdsc = 0
+ cdscb = 0 cdscd = 0 pclm = 0.653425
+ wpclm = -2.221987E-6 pdiblc1 = 0.21098 pdiblc2 = 2E-4
+ pdiblcb = -0.26831 drout = 0.36075 pscbe1 = 9.3731E8
+ pscbe2 = 1.68E-6 pvag = 1.99 delta = 0.0246
+ fprout = 10.125 pdits = 0 pditsl = 0
+ pditsd = 0 lambda = 0 vtl = 0
+ lc = 5E-9 xn = 3 alpha0 = 2.378922E-5
+ walpha0 = -6.485754E-11 alpha1 = 0 beta0 = 26.68934
+ wbeta0 = -1.871056E-5 aigbacc = 1 bigbacc = 0
+ cigbacc = 0 nigbacc = 1 aigbinv = 0.35
+ bigbinv = 0.03 cigbinv = 6E-3 eigbinv = 1.1
+ nigbinv = 3 aigc = 0.43 bigc = 0.054
+ cigc = 0.075 aigsd = 0.43 bigsd = 0.054
+ cigsd = 0.075 dlcig = 0 nigc = 1
+ poxedge = 1 pigcd = 1 ntox = 1
+ toxref = 1.16E-8 agidl = 5.06E-11 bgidl = 1.058E9
+ cgidl = 4E3 egidl = 0.8 noia = 2.6E41
+ noib = 0 noic = 0 em = 4.1E7
+ af = 1 ef = 0.89 kf = 0
+ lintnoi = 0 tnoia = 7.5E6 tnoib = 7.2E6
+ ntnoi = 1 rnoia = 0.794 rnoib = 0.38
+ xpart = 0 cgso = {2.754679E-10/sw_func_tox_hv_ratio} cgdo = {2.754679E-10/sw_func_tox_hv_ratio}
+ cgbo = {0/sw_func_tox_hv_ratio} ckappas = 0.6 cf = 0
+ clc = 1E-7 cle = 0.6 dlc = 6.5995E-8
+ dwc = 0 vfbcv = -1 noff = 4
+ voffcv = -0.4104 acde = 0.4176 moin = 15
+ cgsl = {4.49025E-11/sw_func_tox_hv_ratio} cgdl = {4.49025E-11/sw_func_tox_hv_ratio} ijthsrev = 0.1
+ ijthsfwd = 0.1 xjbvs = 1 bvs = 12.636
+ jss = 3.75E-4 jsws = 5.84E-11 cjs = {8.310E-04*sw_func_nsd_pw_cj}
+ mjs = 0.295 mjsws = 0.037586 cjsws = {8.643094E-11*sw_func_nsd_pw_cj}
+ cjswgs = {5.47776E-11*sw_func_nsd_pw_cj} mjswgs = 0.78692 pbs = 0.72468
+ pbsws = 0.29067 pbswgs = 0.54958 xrcrg1 = 12
+ xrcrg2 = 1 rbpb = 50 rbpd = 50
+ rbps = 50 rbdb = 50 rbsb = 50
+ gbmin = 1E-12 tnom = 30 ute = -1.2986
+ kt1 = -0.40273 kt1l = 0 kt2 = -0.019151
+ ua1 = 3.0044E-9 ub1 = -3.7525E-18 uc1 = -5.9821E-11
+ at = 1.798292E5 wat = -0.137958 prt = 0
+ njs = 1.0773 xtis = 0.76 tpb = 1.344E-3
+ tpbsw = 9.9005E-4 tpbswg = 0 tcj = 6.7434E-4
+ tcjsw = 2.493E-4 tcjswg = 0 tvoff = 0
+ tvfbsdoff = 0 saref = 3E-6 sbref = 3E-6
+ wlod = 0 ku0 = -4.5E-8 kvsat = 0.3
+ kvth0 = 1.1E-8 tku0 = 0 llodku0 = 0
+ wlodku0 = 1 llodvth = 0 wlodvth = 1
+ lku0 = 0 wku0 = 2E-7 pku0 = 0
+ lkvth0 = 0 wkvth0 = 6.5E-7 pkvth0 = 0
+ stk2 = 0 lodk2 = 1 steta0 = 0
+ lodeta0 = 1

.model nhv_model.23 nmos
+ level = 54 lmin = 4E-6 lmax = 8E-6 wmin = 5E-6
+ wmax = 7E-6 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 1.16E-8
+ toxm = 1.16E-8 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 1E23 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {2.1346E-8+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {7.6507E-8-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = -4.1292E-9 dwb = -1.6944E-9 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = 0.762108 lvth0 = 9.277268E-8
+ wvth0 = 1.479046E-7 pvth0 = -3.477419E-13 k1 = 0.88325
+ k2 = -3.97195E-2 lk2 = 5.605426E-9 wk2 = -8.91979E-9
+ pk2 = 3.386319E-14 k3 = -0.884 k3b = 0.43
+ w0 = 0 lpe0 = 2.5E-8 lpeb = -2.182E-7
+ vbm = -3 dvtp0 = 0 dvtp1 = 0
+ dvt0 = 0 dvt1 = 0.53 dvt2 = -0.19251
+ dvt0w = 0.16 dvt1w = 6.9091E6 dvt2w = -0.036016
+ vfbsdoff = 0 u0 = 4.01955E-2 lu0 = 8.623308E-9
+ wu0 = 9.474366E-9 pu0 = -2.991986E-14 ua = -5.25742E-10
+ lua = 1.162239E-15 wua = 2.950861E-15 pua = -5.773427E-21
+ ub = 2.320551E-18 lub = -1.30522E-24 wub = -3.953067E-24
+ pub = 7.134436E-30 uc = 6.6204E-11 ud = 0
+ up = 0 lp = 1 eu = 1.67
+ vsat = 1.422156E5 lvsat = -0.18046 wvsat = -0.220873
+ pvsat = 9.929907E-7 a0 = 1.540926 la0 = -2.440438E-6
+ wa0 = -3.529545E-6 pa0 = 1.201016E-11 ags = 0.202417
+ lags = -2.552557E-7 wags = -3.503067E-7 pags = 1.631303E-12
+ b0 = 3.2933E-8 b1 = 0 keta = -2.934507E-3
+ lketa = -1.106028E-7 wketa = -9.972365E-8 pketa = 5.482922E-13
+ a1 = 0 a2 = 0.659726 rdsw = 724.62
+ rdswmin = 0 rdw = 0 rdwmin = 0
+ rsw = 0 rswmin = 0 prwb = 0.05626
+ prwg = 0.048 wr = 1 voff = -0.20613
+ voffl = -4.257949E-7 minv = 0 nfactor = 0.928619
+ lnfactor = -1.546104E-7 wnfactor = 5.807447E-7 pnfactor = -1.47452E-12
+ eta0 = 0.032 etab = -0.01932 dsub = 0.504
+ cit = -8E-4 cdsc = 0 cdscb = 0
+ cdscd = 0 pclm = 0.395514 lpclm = 2.023824E-6
+ wpclm = -9.434429E-7 ppclm = -1.003272E-11 pdiblc1 = 0.21098
+ pdiblc2 = 2E-4 pdiblcb = -0.26831 drout = 0.36075
+ pscbe1 = 9.3731E8 pscbe2 = 1.68E-6 pvag = 1.99
+ delta = 0.0246 fprout = 10.125 pdits = 0
+ pditsl = 0 pditsd = 0 lambda = 0
+ vtl = 0 lc = 5E-9 xn = 3
+ alpha0 = 3.551293E-5 lalpha0 = -9.199578E-11 walpha0 = -1.46423E-10
+ palpha0 = 6.40043E-16 alpha1 = 0 beta0 = 26.801484
+ lbeta0 = -8.799943E-7 wbeta0 = -3.688782E-5 pbeta0 = 1.426367E-10
+ aigbacc = 1 bigbacc = 0 cigbacc = 0
+ nigbacc = 1 aigbinv = 0.35 bigbinv = 0.03
+ cigbinv = 6E-3 eigbinv = 1.1 nigbinv = 3
+ aigc = 0.43 bigc = 0.054 cigc = 0.075
+ aigsd = 0.43 bigsd = 0.054 cigsd = 0.075
+ dlcig = 0 nigc = 1 poxedge = 1
+ pigcd = 1 ntox = 1 toxref = 1.16E-8
+ agidl = 5.06E-11 bgidl = 1.058E9 cgidl = 4E3
+ egidl = 0.8 noia = 2.6E41 noib = 0
+ noic = 0 em = 4.1E7 af = 1
+ ef = 0.89 kf = 0 lintnoi = 0
+ tnoia = 7.5E6 tnoib = 7.2E6 ntnoi = 1
+ rnoia = 0.794 rnoib = 0.38 xpart = 0
+ cgso = {2.754679E-10/sw_func_tox_hv_ratio} cgdo = {2.754679E-10/sw_func_tox_hv_ratio} cgbo = {0/sw_func_tox_hv_ratio}
+ ckappas = 0.6 cf = 0 clc = 1E-7
+ cle = 0.6 dlc = 6.5995E-8 dwc = 0
+ vfbcv = -1 noff = 4 voffcv = -0.4104
+ acde = 0.4176 moin = 15 cgsl = {4.49025E-11/sw_func_tox_hv_ratio}
+ cgdl = {4.49025E-11/sw_func_tox_hv_ratio} ijthsrev = 0.1 ijthsfwd = 0.1
+ xjbvs = 1 bvs = 12.636 jss = 3.75E-4
+ jsws = 5.84E-11 cjs = {8.310E-04*sw_func_nsd_pw_cj} mjs = 0.295
+ mjsws = 0.037586 cjsws = {8.643094E-11*sw_func_nsd_pw_cj} cjswgs = {5.47776E-11*sw_func_nsd_pw_cj}
+ mjswgs = 0.78692 pbs = 0.72468 pbsws = 0.29067
+ pbswgs = 0.54958 xrcrg1 = 12 xrcrg2 = 1
+ rbpb = 50 rbpd = 50 rbps = 50
+ rbdb = 50 rbsb = 50 gbmin = 1E-12
+ tnom = 30 ute = -1.33707 lute = 3.018725E-7
+ kt1 = -0.414271 lkt1 = 9.056174E-8 kt1l = 0
+ kt2 = -0.019151 ua1 = 3.0044E-9 ub1 = -3.7525E-18
+ uc1 = -5.9821E-11 at = 2.758396E5 lat = -0.753392
+ wat = -0.270639 pat = 1.041144E-6 prt = 0
+ njs = 1.0773 xtis = 0.76 tpb = 1.344E-3
+ tpbsw = 9.9005E-4 tpbswg = 0 tcj = 6.7434E-4
+ tcjsw = 2.493E-4 tcjswg = 0 tvoff = 0
+ tvfbsdoff = 0 saref = 3E-6 sbref = 3E-6
+ wlod = 0 ku0 = -4.5E-8 kvsat = 0.3
+ kvth0 = 1.1E-8 tku0 = 0 llodku0 = 0
+ wlodku0 = 1 llodvth = 0 wlodvth = 1
+ lku0 = 0 wku0 = 2E-7 pku0 = 0
+ lkvth0 = 0 wkvth0 = 6.5E-7 pkvth0 = 0
+ stk2 = 0 lodk2 = 1 steta0 = 0
+ lodeta0 = 1

.model nhv_model.24 nmos
+ level = 54 lmin = 2E-6 lmax = 4E-6 wmin = 5E-6
+ wmax = 7E-6 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 1.16E-8
+ toxm = 1.16E-8 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 1E23 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {2.1346E-8+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {7.6507E-8-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = -4.1292E-9 dwb = -1.6944E-9 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = 0.794536 lvth0 = -3.197647E-8
+ wvth0 = 3.266763E-8 pvth0 = 9.557316E-14 k1 = 0.88325
+ k2 = -4.32634E-2 lk2 = 1.923862E-8 wk2 = 4.832354E-9
+ pk2 = -1.904111E-14 k3 = -0.884 k3b = 0.43
+ w0 = 0 lpe0 = 2.5E-8 lpeb = -2.182E-7
+ vbm = -3 dvtp0 = 0 dvtp1 = 0
+ dvt0 = 0 dvt1 = 0.53 dvt2 = -0.19251
+ dvt0w = 0.16 dvt1w = 6.9091E6 dvt2w = -0.036016
+ vfbsdoff = 0 u0 = 4.38512E-2 lu0 = -5.440143E-9
+ wu0 = -7.565337E-9 pu0 = 3.563163E-14 ua = 1.215733E-10
+ lua = -1.327973E-15 wua = -1.08392E-16 pua = 5.995476E-21
+ ub = 1.558319E-18 lub = 1.627077E-24 wub = -6.00617E-26
+ pub = -7.8419E-30 uc = 6.6204E-11 ud = 0
+ up = 0 lp = 1 eu = 1.67
+ vsat = 7.304387E4 lvsat = 8.56425E-2 wvsat = 0.144267
+ pvsat = -4.116998E-7 a0 = 0.277443 la0 = 2.420165E-6
+ wa0 = 1.385138E-6 pa0 = -6.896553E-12 ags = 0.114213
+ lags = 8.406631E-8 wags = 3.633311E-8 pags = 1.43905E-13
+ b0 = 3.2933E-8 b1 = 0 keta = -5.11015E-2
+ lketa = 7.469484E-8 wketa = 8.232837E-8 pketa = -1.520593E-13
+ a1 = 0 a2 = 0.659726 rdsw = 724.62
+ rdswmin = 0 rdw = 0 rdwmin = 0
+ rsw = 0 rswmin = 0 prwb = 0.05626
+ prwg = 0.048 wr = 1 voff = -0.20613
+ voffl = -4.257949E-7 minv = 0 nfactor = 0.943206
+ lnfactor = -2.107241E-7 wnfactor = 1.261066E-7 pnfactor = 2.744665E-13
+ eta0 = 0.032 etab = -0.01932 dsub = 0.504
+ cit = -8E-4 cdsc = 0 cdscb = 0
+ cdscd = 0 pclm = 1.58199 lpclm = -2.540535E-6
+ wpclm = -6.825173E-6 ppclm = 1.259421E-11 pdiblc1 = 0.21098
+ pdiblc2 = 2E-4 pdiblcb = -0.26831 drout = 0.36075
+ pscbe1 = 9.3731E8 pscbe2 = 1.68E-6 pvag = 1.99
+ delta = 0.0246 fprout = 10.125 pdits = 0
+ pditsl = 0 pditsd = 0 lambda = 0
+ vtl = 0 lc = 5E-9 xn = 3
+ alpha0 = 8.950802E-6 lalpha0 = 1.018834E-11 walpha0 = 3.837789E-11
+ palpha0 = -7.088343E-17 alpha1 = 0 beta0 = 23.806628
+ lbeta0 = 1.064117E-5 wbeta0 = 3.648719E-7 pbeta0 = -6.739133E-13
+ aigbacc = 1 bigbacc = 0 cigbacc = 0
+ nigbacc = 1 aigbinv = 0.35 bigbinv = 0.03
+ cigbinv = 6E-3 eigbinv = 1.1 nigbinv = 3
+ aigc = 0.43 bigc = 0.054 cigc = 0.075
+ aigsd = 0.43 bigsd = 0.054 cigsd = 0.075
+ dlcig = 0 nigc = 1 poxedge = 1
+ pigcd = 1 ntox = 1 toxref = 1.16E-8
+ agidl = 5.06E-11 bgidl = 1.058E9 cgidl = 4E3
+ egidl = 0.8 noia = 2.6E41 noib = 0
+ noic = 0 em = 4.1E7 af = 1
+ ef = 0.89 kf = 0 lintnoi = 0
+ tnoia = 7.5E6 tnoib = 7.2E6 ntnoi = 1
+ rnoia = 0.794 rnoib = 0.38 xpart = 0
+ cgso = {2.754679E-10/sw_func_tox_hv_ratio} cgdo = {2.754679E-10/sw_func_tox_hv_ratio} cgbo = {0/sw_func_tox_hv_ratio}
+ ckappas = 0.6 cf = 0 clc = 1E-7
+ cle = 0.6 dlc = 6.5995E-8 dwc = 0
+ vfbcv = -1 noff = 4 voffcv = -0.4104
+ acde = 0.4176 moin = 15 cgsl = {4.49025E-11/sw_func_tox_hv_ratio}
+ cgdl = {4.49025E-11/sw_func_tox_hv_ratio} ijthsrev = 0.1 ijthsfwd = 0.1
+ xjbvs = 1 bvs = 12.636 jss = 3.75E-4
+ jsws = 5.84E-11 cjs = {8.310E-04*sw_func_nsd_pw_cj} mjs = 0.295
+ mjsws = 0.037586 cjsws = {8.643094E-11*sw_func_nsd_pw_cj} cjswgs = {5.47776E-11*sw_func_nsd_pw_cj}
+ mjswgs = 0.78692 pbs = 0.72468 pbsws = 0.29067
+ pbswgs = 0.54958 xrcrg1 = 12 xrcrg2 = 1
+ rbpb = 50 rbpd = 50 rbps = 50
+ rbdb = 50 rbsb = 50 gbmin = 1E-12
+ tnom = 30 ute = -1.22166 lute = -1.421066E-7
+ kt1 = -0.407353 lkt1 = 6.394796E-8 kt1l = 0
+ kt2 = -0.019151 ua1 = 3.0044E-9 ub1 = -3.7525E-18
+ uc1 = -5.9821E-11 at = 1.482596E5 lat = -0.262594
+ wat = -6.37017E-2 pat = 2.450594E-7 prt = 0
+ njs = 1.0773 xtis = 0.76 tpb = 1.344E-3
+ tpbsw = 9.9005E-4 tpbswg = 0 tcj = 6.7434E-4
+ tcjsw = 2.493E-4 tcjswg = 0 tvoff = 0
+ tvfbsdoff = 0 saref = 3E-6 sbref = 3E-6
+ wlod = 0 ku0 = -4.5E-8 kvsat = 0.3
+ kvth0 = 1.1E-8 tku0 = 0 llodku0 = 0
+ wlodku0 = 1 llodvth = 0 wlodvth = 1
+ lku0 = 0 wku0 = 2E-7 pku0 = 0
+ lkvth0 = 0 wkvth0 = 6.5E-7 pkvth0 = 0
+ stk2 = 0 lodk2 = 1 steta0 = 0
+ lodeta0 = 1

.model nhv_model.25 nmos
+ level = 54 lmin = 1E-6 lmax = 2E-6 wmin = 5E-6
+ wmax = 7E-6 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 1.16E-8
+ toxm = 1.16E-8 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 1E23 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {2.1346E-8+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {7.6507E-8-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = -4.1292E-9 dwb = -1.6944E-9 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = 0.751772 lvth0 = 4.700719E-8
+ wvth0 = 2.105803E-7 pvth0 = -2.330291E-13 k1 = 0.88325
+ k2 = -0.061201 lk2 = 5.23691E-8 wk2 = 1.350817E-7
+ pk2 = -2.596097E-13 k3 = -0.884 k3b = 0.43
+ w0 = 0 lpe0 = 2.5E-8 lpeb = -2.182E-7
+ vbm = -3 dvtp0 = 0 dvtp1 = 0
+ dvt0 = 0 dvt1 = 0.53 dvt2 = -0.19251
+ dvt0w = 0.16 dvt1w = 6.9091E6 dvt2w = -0.036016
+ vfbsdoff = 0 u0 = 3.74512E-2 lu0 = 6.380635E-9
+ wu0 = 2.885205E-8 pu0 = -3.163077E-14 ua = -5.907914E-10
+ lua = -1.224592E-17 wua = 3.104826E-15 pua = 6.070681E-23
+ ub = 2.447652E-18 lub = -1.550943E-26 wub = -4.347471E-24
+ pub = 7.688504E-32 uc = 6.6204E-11 ud = 0
+ up = 0 lp = 1 eu = 1.67
+ vsat = 1.390944E5 lvsat = -3.63519E-2 wvsat = -0.176205
+ pvsat = 1.802077E-7 a0 = 1.583728 la0 = 7.474458E-9
+ wa0 = -2.328751E-6 pa0 = -3.705319E-14 ags = 0.190305
+ lags = -5.647556E-8 wags = -3.73338E-8 pags = 2.799667E-13
+ b0 = 3.2933E-8 b1 = 0 keta = -0.01066
+ a1 = 0 a2 = 0.659726 rdsw = 724.62
+ rdswmin = 0 rdw = 0 rdwmin = 0
+ rsw = 0 rswmin = 0 prwb = 0.05626
+ prwg = 0.048 wr = 1 voff = -0.20613
+ voffl = -4.257949E-7 minv = 0 nfactor = 0.952509
+ lnfactor = -2.27907E-7 wnfactor = -3.369932E-7 pnfactor = 1.129805E-12
+ eta0 = 0.032 etab = -0.01932 dsub = 0.504
+ cit = -8E-4 cdsc = 0 cdscb = 0
+ cdscd = 0 pclm = -1.307712 lpclm = 2.796705E-6
+ wpclm = 7.499971E-6 ppclm = -1.386413E-11 pdiblc1 = 0.21098
+ pdiblc2 = 2E-4 pdiblcb = -0.26831 drout = 0.36075
+ pscbe1 = 9.3731E8 pscbe2 = 1.68E-6 pvag = 1.99
+ delta = 0.0246 fprout = 10.125 pdits = 0
+ pditsl = 0 pditsd = 0 lambda = 0
+ vtl = 0 lc = 5E-9 xn = 3
+ alpha0 = 1.787595E-5 lalpha0 = -6.296286E-12 walpha0 = -1.689922E-11
+ palpha0 = 3.121263E-17 alpha1 = 0 beta0 = 20.045328
+ lbeta0 = 1.758824E-5 wbeta0 = 4.720682E-5 pbeta0 = -8.719033E-11
+ aigbacc = 1 bigbacc = 0 cigbacc = 0
+ nigbacc = 1 aigbinv = 0.35 bigbinv = 0.03
+ cigbinv = 6E-3 eigbinv = 1.1 nigbinv = 3
+ aigc = 0.43 bigc = 0.054 cigc = 0.075
+ aigsd = 0.43 bigsd = 0.054 cigsd = 0.075
+ dlcig = 0 nigc = 1 poxedge = 1
+ pigcd = 1 ntox = 1 toxref = 1.16E-8
+ agidl = 5.06E-11 bgidl = 1.058E9 cgidl = 4E3
+ egidl = 0.8 noia = 2.6E41 noib = 0
+ noic = 0 em = 4.1E7 af = 1
+ ef = 0.89 kf = 0 lintnoi = 0
+ tnoia = 7.5E6 tnoib = 7.2E6 ntnoi = 1
+ rnoia = 0.794 rnoib = 0.38 xpart = 0
+ cgso = {2.754679E-10/sw_func_tox_hv_ratio} cgdo = {2.754679E-10/sw_func_tox_hv_ratio} cgbo = {0/sw_func_tox_hv_ratio}
+ ckappas = 0.6 cf = 0 clc = 1E-7
+ cle = 0.6 dlc = 6.5995E-8 dwc = 0
+ vfbcv = -1 noff = 4 voffcv = -0.4104
+ acde = 0.4176 moin = 15 cgsl = {4.49025E-11/sw_func_tox_hv_ratio}
+ cgdl = {4.49025E-11/sw_func_tox_hv_ratio} ijthsrev = 0.1 ijthsfwd = 0.1
+ xjbvs = 1 bvs = 12.636 jss = 3.75E-4
+ jsws = 5.84E-11 cjs = {8.310E-04*sw_func_nsd_pw_cj} mjs = 0.295
+ mjsws = 0.037586 cjsws = {8.643094E-11*sw_func_nsd_pw_cj} cjswgs = {5.47776E-11*sw_func_nsd_pw_cj}
+ mjswgs = 0.78692 pbs = 0.72468 pbsws = 0.29067
+ pbswgs = 0.54958 xrcrg1 = 12 xrcrg2 = 1
+ rbpb = 50 rbpd = 50 rbps = 50
+ rbdb = 50 rbsb = 50 gbmin = 1E-12
+ tnom = 30 ute = -1.2986 kt1 = -0.37273
+ kt1l = 0 kt2 = -0.019151 ua1 = 3.0044E-9
+ ub1 = -3.7525E-18 uc1 = -5.9821E-11 at = -1.748559E4
+ lat = 4.35353E-2 wat = 0.185828 pat = -2.158177E-7
+ prt = 0 njs = 1.0773 xtis = 0.76
+ tpb = 1.344E-3 tpbsw = 9.9005E-4 tpbswg = 0
+ tcj = 6.7434E-4 tcjsw = 2.493E-4 tcjswg = 0
+ tvoff = 0 tvfbsdoff = 0 saref = 3E-6
+ sbref = 3E-6 wlod = 0 ku0 = -4.5E-8
+ kvsat = 0.3 kvth0 = 1.1E-8 tku0 = 0
+ llodku0 = 0 wlodku0 = 1 llodvth = 0
+ wlodvth = 1 lku0 = 0 wku0 = 2E-7
+ pku0 = 0 lkvth0 = 0 wkvth0 = 6.5E-7
+ pkvth0 = 0 stk2 = 0 lodk2 = 1
+ steta0 = 0 lodeta0 = 1

.model nhv_model.26 nmos
+ level = 54 lmin = 8E-7 lmax = 1E-6 wmin = 5E-6
+ wmax = 7E-6 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 1.16E-8
+ toxm = 1.16E-8 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 1E23 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {2.1346E-8+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {7.6507E-8-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = -4.1292E-9 dwb = -1.6944E-9 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = 0.802565 lvth0 = 3.986799E-9
+ wvth0 = -2.215278E-7 pvth0 = 1.329604E-13 k1 = 0.88325
+ k2 = -4.964979E-3 lk2 = 4.737981E-9 wk2 = -1.792105E-7
+ pk2 = 6.591321E-15 k3 = -0.884 k3b = 0.43
+ w0 = 0 lpe0 = 2.5E-8 lpeb = -2.182E-7
+ vbm = -3 dvtp0 = 0 dvtp1 = 0
+ dvt0 = 0 dvt1 = 0.53 dvt2 = -0.19251
+ dvt0w = 0.16 dvt1w = 6.9091E6 dvt2w = -0.036016
+ vfbsdoff = 0 u0 = 8.51559E-2 lu0 = -3.402456E-8
+ wu0 = -2.901043E-7 pu0 = 2.385208E-13 ua = -2.090784E-9
+ lua = 1.258227E-15 wua = 1.350136E-14 pua = -8.74501E-21
+ ub = 1.146453E-17 lub = -7.65268E-24 wub = -7.069064E-23
+ pub = 5.626862E-29 uc = 6.6204E-11 ud = 0
+ up = 0 lp = 1 eu = 1.67
+ vsat = 1.636616E5 lvsat = -0.05716 wvsat = -0.333578
+ pvsat = 3.135012E-7 a0 = 3.11411 la0 = -1.288738E-6
+ wa0 = -1.004736E-5 pa0 = 6.500503E-12 ags = 5.153286E-3
+ lags = 1.003454E-7 wags = 1.241728E-6 pags = -8.033804E-13
+ b0 = 3.2933E-8 b1 = 0 keta = -0.01066
+ a1 = 0 a2 = 0.659726 rdsw = 724.62
+ rdswmin = 0 rdw = 0 rdwmin = 0
+ rsw = 0 rswmin = 0 prwb = 0.05626
+ prwg = 0.048 wr = 1 voff = -0.20613
+ voffl = -4.257949E-7 minv = 0 nfactor = 7.72381E-2
+ lnfactor = 5.134352E-7 wnfactor = 5.324208E-6 pnfactor = -3.665152E-12
+ eta0 = 0.032 etab = -0.01932 dsub = 0.504
+ cit = -8E-4 cdsc = 0 cdscb = 0
+ cdscd = 0 pclm = 7.181289 lpclm = -4.39336E-6
+ wpclm = -5.189567E-5 ppclm = 3.644315E-11 pdiblc1 = 0.21098
+ pdiblc2 = 2E-4 pdiblcb = -0.26831 drout = 0.36075
+ pscbe1 = 9.3731E8 pscbe2 = 1.68E-6 pvag = 1.99
+ delta = 0.0246 fprout = 10.125 pdits = 0
+ pditsl = 0 pditsd = 0 lambda = 0
+ vtl = 0 lc = 5E-9 xn = 3
+ alpha0 = -3.513327E-5 lalpha0 = 3.860178E-11 walpha0 = 2.458838E-10
+ palpha0 = -1.913609E-16 alpha1 = 0 beta0 = 69.900989
+ lbeta0 = -2.463881E-5 wbeta0 = -3.184852E-4 pbeta0 = 2.225457E-10
+ aigbacc = 1 bigbacc = 0 cigbacc = 0
+ nigbacc = 1 aigbinv = 0.35 bigbinv = 0.03
+ cigbinv = 6E-3 eigbinv = 1.1 nigbinv = 3
+ aigc = 0.43 bigc = 0.054 cigc = 0.075
+ aigsd = 0.43 bigsd = 0.054 cigsd = 0.075
+ dlcig = 0 nigc = 1 poxedge = 1
+ pigcd = 1 ntox = 1 toxref = 1.16E-8
+ agidl = 5.06E-11 bgidl = 1.058E9 cgidl = 4E3
+ egidl = 0.8 noia = 2.6E41 noib = 0
+ noic = 0 em = 4.1E7 af = 1
+ ef = 0.89 kf = 0 lintnoi = 0
+ tnoia = 7.5E6 tnoib = 7.2E6 ntnoi = 1
+ rnoia = 0.794 rnoib = 0.38 xpart = 0
+ cgso = {2.754679E-10/sw_func_tox_hv_ratio} cgdo = {2.754679E-10/sw_func_tox_hv_ratio} cgbo = {0/sw_func_tox_hv_ratio}
+ ckappas = 0.6 cf = 0 clc = 1E-7
+ cle = 0.6 dlc = 6.5995E-8 dwc = 0
+ vfbcv = -1 noff = 4 voffcv = -0.4104
+ acde = 0.4176 moin = 15 cgsl = {4.49025E-11/sw_func_tox_hv_ratio}
+ cgdl = {4.49025E-11/sw_func_tox_hv_ratio} ijthsrev = 0.1 ijthsfwd = 0.1
+ xjbvs = 1 bvs = 12.636 jss = 3.75E-4
+ jsws = 5.84E-11 cjs = {8.310E-04*sw_func_nsd_pw_cj} mjs = 0.295
+ mjsws = 0.037586 cjsws = {8.643094E-11*sw_func_nsd_pw_cj} cjswgs = {5.47776E-11*sw_func_nsd_pw_cj}
+ mjswgs = 0.78692 pbs = 0.72468 pbsws = 0.29067
+ pbswgs = 0.54958 xrcrg1 = 12 xrcrg2 = 1
+ rbpb = 50 rbpd = 50 rbps = 50
+ rbdb = 50 rbsb = 50 gbmin = 1E-12
+ tnom = 30 ute = -1.87814 lute = 4.908622E-7
+ wute = 2.872958E-6 pute = -2.433355E-12 kt1 = -0.218834
+ lkt1 = -1.303474E-7 wkt1 = -1.115712E-6 pkt1 = 9.449923E-13
+ kt1l = 0 kt2 = -0.019151 ua1 = 1.417545E-8
+ lua1 = -9.461726E-15 wua1 = -5.537835E-14 pua1 = 4.690469E-20
+ ub1 = -2.80931E-17 lub1 = 2.061615E-23 wub1 = 1.174566E-22
+ pub1 = -9.948406E-29 uc1 = -5.9821E-11 at = 2.149895E5
+ lat = -0.153368 wat = -1.441305 pat = 1.16234E-6
+ prt = 0 njs = 1.0773 xtis = 0.76
+ tpb = 1.344E-3 tpbsw = 9.9005E-4 tpbswg = 0
+ tcj = 6.7434E-4 tcjsw = 2.493E-4 tcjswg = 0
+ tvoff = 0 tvfbsdoff = 0 saref = 3E-6
+ sbref = 3E-6 wlod = 0 ku0 = -4.5E-8
+ kvsat = 0.3 kvth0 = 1.1E-8 tku0 = 0
+ llodku0 = 0 wlodku0 = 1 llodvth = 0
+ wlodvth = 1 lku0 = 0 wku0 = 2E-7
+ pku0 = 0 lkvth0 = 0 wkvth0 = 6.5E-7
+ pkvth0 = 0 stk2 = 0 lodk2 = 1
+ steta0 = 0 lodeta0 = 1

.model nhv_model.27 nmos
+ level = 54 lmin = 6E-7 lmax = 8E-7 wmin = 5E-6
+ wmax = 7E-6 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 1.16E-8
+ toxm = 1.16E-8 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 1E23 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {2.1346E-8+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {7.6507E-8-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = -4.1292E-9 dwb = -1.6944E-9 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = 0.808727 wvth0 = -1.602038E-8
+ k1 = 0.88325 k2 = 2.358179E-3 wk2 = -1.690228E-7
+ k3 = -0.884 k3b = 0.43 w0 = 0
+ lpe0 = 2.5E-8 lpeb = -2.182E-7 vbm = -3
+ dvtp0 = 0 dvtp1 = 0 dvt0 = 0
+ dvt1 = 0.53 dvt2 = -0.19251 dvt0w = 0.16
+ dvt1w = 6.9091E6 dvt2w = -0.036016 vfbsdoff = 0
+ u0 = 3.25665E-2 wu0 = 7.856023E-8 ua = -1.460326E-10
+ wua = -1.517884E-17 ub = -3.636685E-19 wub = 1.627974E-23
+ uc = 6.6204E-11 ud = 0 up = 0
+ lp = 1 eu = 1.67 vsat = 7.531348E4
+ wvsat = 0.150978 a0 = 1.1222 ags = 0.16025
+ b0 = 3.2933E-8 b1 = 0 keta = -0.01066
+ a1 = 0 a2 = 0.659726 rdsw = 724.62
+ rdswmin = 0 rdw = 0 rdwmin = 0
+ rsw = 0 rswmin = 0 prwb = 0.05626
+ prwg = 0.048 wr = 1 voff = -0.20613
+ voffl = -4.257949E-7 minv = 0 nfactor = 0.870818
+ wnfactor = -3.407564E-7 eta0 = 0.032 etab = -0.01932
+ dsub = 0.504 cit = -8E-4 cdsc = 0
+ cdscb = 0 cdscd = 0 pclm = 0.390786
+ wpclm = 4.431903E-6 pdiblc1 = 0.21098 pdiblc2 = 2E-4
+ pdiblcb = -0.26831 drout = 0.36075 pscbe1 = 9.3731E8
+ pscbe2 = 1.68E-6 pvag = 1.99 delta = 0.0246
+ fprout = 10.125 pdits = 0 pditsl = 0
+ pditsd = 0 lambda = 0 vtl = 0
+ lc = 5E-9 xn = 3 alpha0 = 2.453075E-5
+ walpha0 = -4.988909E-11 alpha1 = 0 beta0 = 31.818549
+ wbeta0 = 2.548775E-5 aigbacc = 1 bigbacc = 0
+ cigbacc = 0 nigbacc = 1 aigbinv = 0.35
+ bigbinv = 0.03 cigbinv = 6E-3 eigbinv = 1.1
+ nigbinv = 3 aigc = 0.43 bigc = 0.054
+ cigc = 0.075 aigsd = 0.43 bigsd = 0.054
+ cigsd = 0.075 dlcig = 0 nigc = 1
+ poxedge = 1 pigcd = 1 ntox = 1
+ toxref = 1.16E-8 agidl = 5.06E-11 bgidl = 1.058E9
+ cgidl = 4E3 egidl = 0.8 noia = 2.6E41
+ noib = 0 noic = 0 em = 4.1E7
+ af = 1 ef = 0.89 kf = 0
+ lintnoi = 0 tnoia = 7.5E6 tnoib = 7.2E6
+ ntnoi = 1 rnoia = 0.794 rnoib = 0.38
+ xpart = 0 cgso = {2.754679E-10/sw_func_tox_hv_ratio} cgdo = {2.754679E-10/sw_func_tox_hv_ratio}
+ cgbo = {0/sw_func_tox_hv_ratio} ckappas = 0.6 cf = 0
+ clc = 1E-7 cle = 0.6 dlc = 6.5995E-8
+ dwc = 0 vfbcv = -1 noff = 4
+ voffcv = -0.4104 acde = 0.4176 moin = 15
+ cgsl = {4.49025E-11/sw_func_tox_hv_ratio} cgdl = {4.49025E-11/sw_func_tox_hv_ratio} ijthsrev = 0.1
+ ijthsfwd = 0.1 xjbvs = 1 bvs = 12.636
+ jss = 3.75E-4 jsws = 5.84E-11 cjs = {8.310E-04*sw_func_nsd_pw_cj}
+ mjs = 0.295 mjsws = 0.037586 cjsws = {8.643094E-11*sw_func_nsd_pw_cj}
+ cjswgs = {5.47776E-11*sw_func_nsd_pw_cj} mjswgs = 0.78692 pbs = 0.72468
+ pbsws = 0.29067 pbswgs = 0.54958 xrcrg1 = 12
+ xrcrg2 = 1 rbpb = 50 rbpd = 50
+ rbps = 50 rbdb = 50 rbsb = 50
+ gbmin = 1E-12 tnom = 30 ute = -1.119449
+ wute = -8.881051E-7 kt1 = -0.420303 wkt1 = 3.448952E-7
+ kt1l = 0 kt2 = -0.019151 ua1 = -4.488598E-10
+ wua1 = 1.711887E-14 ub1 = 3.771806E-18 wub1 = -3.630884E-23
+ uc1 = -5.9821E-11 at = -2.206027E4 wat = 0.355242
+ prt = 0 njs = 1.0773 xtis = 0.76
+ tpb = 1.344E-3 tpbsw = 9.9005E-4 tpbswg = 0
+ tcj = 6.7434E-4 tcjsw = 2.493E-4 tcjswg = 0
+ tvoff = 0 tvfbsdoff = 0 saref = 1.81E-6
+ sbref = 1.81E-6 wlod = 0 ku0 = -4.5E-8
+ kvsat = 0.3 kvth0 = 1.1E-8 tku0 = 0
+ llodku0 = 0 wlodku0 = 1 llodvth = 0
+ wlodvth = 1 lku0 = 0 wku0 = 2E-7
+ pku0 = 0 lkvth0 = 0 wkvth0 = 6.5E-7
+ pkvth0 = 0 stk2 = 0 lodk2 = 1
+ steta0 = 0 lodeta0 = 1

.model nhv_model.28 nmos
+ level = 54 lmin = 5E-7 lmax = 6E-7 wmin = 5E-6
+ wmax = 7E-6 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 1.16E-8
+ toxm = 1.16E-8 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 1E23 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {2.1346E-8+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {7.6507E-8-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = -4.1292E-9 dwb = -1.6944E-9 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = 0.879689 lvth0 = -3.171908E-8
+ wvth0 = -3.678015E-7 pvth0 = 1.572412E-13 k1 = 0.88325
+ k2 = 0.136907 lk2 = -6.014162E-8 wk2 = -8.360247E-7
+ pk2 = 2.981405E-13 k3 = -0.884 k3b = 0.43
+ w0 = 0 lpe0 = 2.5E-8 lpeb = -2.182E-7
+ vbm = -3 dvtp0 = 0 dvtp1 = 0
+ dvt0 = 0 dvt1 = 0.53 dvt2 = -0.19251
+ dvt0w = 0.16 dvt1w = 6.9091E6 dvt2w = -0.036016
+ vfbsdoff = 0 u0 = -2.99258E-2 lu0 = 2.793318E-8
+ wu0 = 3.883538E-7 pu0 = -1.384734E-13 ua = -1.216409E-10
+ lua = -1.090275E-17 wua = -1.36096E-16 pua = 5.40483E-23
+ ub = -1.223966E-17 lub = 5.3084E-24 wub = 7.515267E-23
+ pub = -2.631537E-29 uc = 6.6204E-11 ud = 0
+ up = 0 lp = 1 eu = 1.67
+ vsat = -1.947075E4 lvsat = 4.23672E-2 wvsat = 0.620853
+ pvsat = -2.100274E-7 a0 = 1.1222 ags = 0.16025
+ b0 = 3.2933E-8 b1 = 0 keta = -0.01066
+ a1 = 0 a2 = 0.659726 rdsw = 724.62
+ rdswmin = 0 rdw = 0 rdwmin = 0
+ rsw = 0 rswmin = 0 prwb = 0.05626
+ prwg = 0.048 wr = 1 voff = -0.20613
+ voffl = -4.257949E-7 minv = 0 nfactor = 1.4846
+ lnfactor = -2.74352E-7 wnfactor = -3.383463E-6 pnfactor = 1.360047E-12
+ eta0 = 0.032 etab = -0.01932 dsub = 0.504
+ cit = -8E-4 cdsc = 0 cdscb = 0
+ cdscd = 0 pclm = -2.711318 lpclm = 1.386597E-6
+ wpclm = 1.980999E-5 ppclm = -6.873788E-12 pdiblc1 = 0.21098
+ pdiblc2 = 2E-4 pdiblcb = -0.26831 drout = 0.36075
+ pscbe1 = 9.3731E8 pscbe2 = 1.68E-6 pvag = 1.99
+ delta = 0.0246 fprout = 10.125 pdits = 0
+ pditsl = 0 pditsd = 0 lambda = 0
+ vtl = 0 lc = 5E-9 xn = 3
+ alpha0 = 5.945054E-5 lalpha0 = -1.560866E-11 walpha0 = -2.229972E-10
+ palpha0 = 7.737692E-17 alpha1 = 0 beta0 = 13.978436
+ lbeta0 = 7.974281E-6 wbeta0 = 1.139267E-4 pbeta0 = -3.953097E-11
+ aigbacc = 1 bigbacc = 0 cigbacc = 0
+ nigbacc = 1 aigbinv = 0.35 bigbinv = 0.03
+ cigbinv = 6E-3 eigbinv = 1.1 nigbinv = 3
+ aigc = 0.43 bigc = 0.054 cigc = 0.075
+ aigsd = 0.43 bigsd = 0.054 cigsd = 0.075
+ dlcig = 0 nigc = 1 poxedge = 1
+ pigcd = 1 ntox = 1 toxref = 1.16E-8
+ agidl = 5.06E-11 bgidl = 1.058E9 cgidl = 4E3
+ egidl = 0.8 noia = 2.6E41 noib = 0
+ noic = 0 em = 4.1E7 af = 1
+ ef = 0.89 kf = 0 lintnoi = 0
+ tnoia = 7.5E6 tnoib = 7.2E6 ntnoi = 1
+ rnoia = 0.794 rnoib = 0.38 xpart = 0
+ cgso = {2.754679E-10/sw_func_tox_hv_ratio} cgdo = {2.754679E-10/sw_func_tox_hv_ratio} cgbo = {0/sw_func_tox_hv_ratio}
+ ckappas = 0.6 cf = 0 clc = 1E-7
+ cle = 0.6 dlc = 6.5995E-8 dwc = 0
+ vfbcv = -1 noff = 4 voffcv = -0.4104
+ acde = 0.4176 moin = 15 cgsl = {4.49025E-11/sw_func_tox_hv_ratio}
+ cgdl = {4.49025E-11/sw_func_tox_hv_ratio} ijthsrev = 0.1 ijthsfwd = 0.1
+ xjbvs = 1 bvs = 12.636 jss = 3.75E-4
+ jsws = 5.84E-11 cjs = {8.310E-04*sw_func_nsd_pw_cj} mjs = 0.295
+ mjsws = 0.037586 cjsws = {8.643094E-11*sw_func_nsd_pw_cj} cjswgs = {5.47776E-11*sw_func_nsd_pw_cj}
+ mjswgs = 0.78692 pbs = 0.72468 pbsws = 0.29067
+ pbswgs = 0.54958 xrcrg1 = 12 xrcrg2 = 1
+ rbpb = 50 rbpd = 50 rbps = 50
+ rbdb = 50 rbsb = 50 gbmin = 1E-12
+ tnom = 30 ute = -0.497822 lute = -2.778589E-7
+ wute = -3.969705E-6 pute = 1.377432E-12 kt1 = -0.661712
+ lkt1 = 1.079064E-7 wkt1 = 1.541633E-6 pkt1 = -5.349251E-13
+ kt1l = 0 kt2 = -0.019151 ua1 = -1.243119E-8
+ lua1 = 5.355933E-15 wua1 = 7.651896E-14 pua1 = -2.655101E-20
+ ub1 = 2.918612E-17 lub1 = -1.135984E-23 wub1 = -1.622954E-22
+ pub1 = 5.631424E-29 uc1 = -5.9821E-11 at = -1.548351E5
+ lat = 5.93485E-2 wat = 1.013448 pat = -2.942088E-7
+ prt = 0 njs = 1.0773 xtis = 0.76
+ tpb = 1.344E-3 tpbsw = 9.9005E-4 tpbswg = 0
+ tcj = 6.7434E-4 tcjsw = 2.493E-4 tcjswg = 0
+ tvoff = 0 tvfbsdoff = 0 saref = 1.81E-6
+ sbref = 1.81E-6 wlod = 0 ku0 = -4.5E-8
+ kvsat = 0.3 kvth0 = 1.1E-8 tku0 = 0
+ llodku0 = 0 wlodku0 = 1 llodvth = 0
+ wlodvth = 1 lku0 = 0 wku0 = 2E-7
+ pku0 = 0 lkvth0 = 0 wkvth0 = 6.5E-7
+ pkvth0 = 0 stk2 = 0 lodk2 = 1
+ steta0 = 0 lodeta0 = 1

.model nhv_model.29 nmos
+ level = 54 lmin = 8E-6 lmax = 2.02E-5 wmin = 3E-6
+ wmax = 5E-6 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 1.16E-8
+ toxm = 1.16E-8 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 1E23 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {2.1346E-8+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {7.6507E-8-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = -4.1292E-9 dwb = -1.6944E-9 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = 0.795471 k1 = 0.88325
+ k2 = -4.22451E-2 wk2 = 1.145701E-8 k3 = -0.884
+ k3b = 0.43 w0 = 0 lpe0 = 2.5E-8
+ lpeb = -2.182E-7 vbm = -3 dvtp0 = 0
+ dvtp1 = 0 dvt0 = 0 dvt1 = 0.53
+ dvt2 = -0.19251 dvt0w = 0.16 dvt1w = 6.9091E6
+ dvt2w = -0.036016 vfbsdoff = 0 u0 = 4.54415E-2
+ wu0 = -1.489654E-8 ua = 3.903403E-10 wua = -1.591951E-15
+ ub = 1.192567E-18 wub = 1.723324E-24 uc = 6.6204E-11
+ ud = 0 up = 0 lp = 1
+ eu = 1.67 vsat = 1.329658E5 wvsat = -0.16248
+ a0 = 0.626333 wa0 = 9.93178E-7 ags = 0.107788
+ wags = 1.654318E-7 b0 = 3.2933E-8 b1 = 0
+ keta = -1.22879E-2 wketa = -5.335611E-8 a1 = 0
+ a2 = 0.659726 rdsw = 724.62 rdswmin = 0
+ rdw = 0 rdwmin = 0 rsw = 0
+ rswmin = 0 prwb = 0.05626 prwg = 0.048
+ wr = 1 voff = -0.20613 voffl = -4.257949E-7
+ minv = 0 nfactor = 0.984478 wnfactor = 1.825206E-8
+ eta0 = 0.032 etab = -0.01932 dsub = 0.504
+ cit = -8E-4 cdsc = 0 cdscb = 0
+ cdscd = 0 pclm = -0.821222 wpclm = 5.088292E-6
+ pdiblc1 = 0.21098 pdiblc2 = 2E-4 pdiblcb = -0.26831
+ drout = 0.36075 pscbe1 = 9.3731E8 pscbe2 = 1.68E-6
+ pvag = 1.99 delta = 0.0246 fprout = 10.125
+ pdits = 0 pditsl = 0 pditsd = 0
+ lambda = 0 vtl = 0 lc = 5E-9
+ xn = 3 alpha0 = 5.144782E-6 walpha0 = 2.756867E-11
+ alpha1 = 0 beta0 = 21.606391 wbeta0 = 6.487177E-6
+ aigbacc = 1 bigbacc = 0 cigbacc = 0
+ nigbacc = 1 aigbinv = 0.35 bigbinv = 0.03
+ cigbinv = 6E-3 eigbinv = 1.1 nigbinv = 3
+ aigc = 0.43 bigc = 0.054 cigc = 0.075
+ aigsd = 0.43 bigsd = 0.054 cigsd = 0.075
+ dlcig = 0 nigc = 1 poxedge = 1
+ pigcd = 1 ntox = 1 toxref = 1.16E-8
+ agidl = 5.06E-11 bgidl = 1.058E9 cgidl = 4E3
+ egidl = 0.8 noia = 2.6E41 noib = 0
+ noic = 0 em = 4.1E7 af = 1
+ ef = 0.89 kf = 0 lintnoi = 0
+ tnoia = 7.5E6 tnoib = 7.2E6 ntnoi = 1
+ rnoia = 0.794 rnoib = 0.38 xpart = 0
+ cgso = {2.754679E-10/sw_func_tox_hv_ratio} cgdo = {2.754679E-10/sw_func_tox_hv_ratio} cgbo = {0/sw_func_tox_hv_ratio}
+ ckappas = 0.6 cf = 0 clc = 1E-7
+ cle = 0.6 dlc = 6.5995E-8 dwc = 0
+ vfbcv = -1 noff = 4 voffcv = -0.4104
+ acde = 0.4176 moin = 15 cgsl = {4.49025E-11/sw_func_tox_hv_ratio}
+ cgdl = {4.49025E-11/sw_func_tox_hv_ratio} ijthsrev = 0.1 ijthsfwd = 0.1
+ xjbvs = 1 bvs = 12.636 jss = 3.75E-4
+ jsws = 5.84E-11 cjs = {8.310E-04*sw_func_nsd_pw_cj} mjs = 0.295
+ mjsws = 0.037586 cjsws = {8.643094E-11*sw_func_nsd_pw_cj} cjswgs = {5.47776E-11*sw_func_nsd_pw_cj}
+ mjswgs = 0.78692 pbs = 0.72468 pbsws = 0.29067
+ pbswgs = 0.54958 xrcrg1 = 12 xrcrg2 = 1
+ rbpb = 50 rbpd = 50 rbps = 50
+ rbdb = 50 rbsb = 50 gbmin = 1E-12
+ tnom = 30 ute = -1.2986 kt1 = -0.40273
+ kt1l = 0 kt2 = -0.019151 ua1 = 3.0044E-9
+ ub1 = -3.7525E-18 uc1 = -5.9821E-11 at = 2.087803E5
+ wat = -0.281478 prt = 0 njs = 1.0773
+ xtis = 0.76 tpb = 1.344E-3 tpbsw = 9.9005E-4
+ tpbswg = 0 tcj = 6.7434E-4 tcjsw = 2.493E-4
+ tcjswg = 0 tvoff = 0 tvfbsdoff = 0
+ saref = 3E-6 sbref = 3E-6 wlod = 0
+ ku0 = -4.5E-8 kvsat = 0.3 kvth0 = 1.1E-8
+ tku0 = 0 llodku0 = 0 wlodku0 = 1
+ llodvth = 0 wlodvth = 1 lku0 = 0
+ wku0 = 2E-7 pku0 = 0 lkvth0 = 0
+ wkvth0 = 6.5E-7 pkvth0 = 0 stk2 = 0
+ lodk2 = 1 steta0 = 0 lodeta0 = 1

.model nhv_model.30 nmos
+ level = 54 lmin = 4E-6 lmax = 8E-6 wmin = 3E-6
+ wmax = 5E-6 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 1.16E-8
+ toxm = 1.16E-8 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 1E23 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {2.1346E-8+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {7.6507E-8-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = -4.1292E-9 dwb = -1.6944E-9 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = 0.79091 lvth0 = 2.326141E-8
+ wvth0 = 5.122447E-9 pvth0 = -3.153195E-15 k1 = 0.88325
+ k2 = -4.37346E-2 lk2 = 1.168761E-8 wk2 = 1.098398E-8
+ pk2 = 3.711919E-15 k3 = -0.884 k3b = 0.43
+ w0 = 0 lpe0 = 2.5E-8 lpeb = -2.182E-7
+ vbm = -3 dvtp0 = 0 dvtp1 = 0
+ dvt0 = 0 dvt1 = 0.53 dvt2 = -0.19251
+ dvt0w = 0.16 dvt1w = 6.9091E6 dvt2w = -0.036016
+ vfbsdoff = 0 u0 = 4.47425E-2 lu0 = 5.48471E-9
+ wu0 = -1.306642E-8 pu0 = -1.436087E-14 ua = 3.91171E-10
+ lua = -6.518951E-18 wua = -1.594559E-15 pua = 2.046811E-23
+ ub = 1.165416E-18 lub = 2.130518E-25 wub = 1.773293E-24
+ pub = -3.921025E-31 uc = 6.6204E-11 ud = 0
+ up = 0 lp = 1 eu = 1.67
+ vsat = 1.381186E5 lvsat = -4.04335E-2 wvsat = -0.200563
+ pvsat = 2.988344E-7 a0 = 0.628541 la0 = -1.732636E-8
+ wa0 = 9.934261E-7 pa0 = -1.947236E-15 ags = 0.101061
+ lags = 5.278859E-8 wags = 1.521487E-7 pags = 1.042325E-13
+ b0 = 3.2933E-8 b1 = 0 keta = -1.22879E-2
+ wketa = -5.335611E-8 a1 = 0 a2 = 0.659726
+ rdsw = 724.62 rdswmin = 0 rdw = 0
+ rdwmin = 0 rsw = 0 rswmin = 0
+ prwb = 0.05626 prwg = 0.048 wr = 1
+ voff = -0.20613 voffl = -4.257949E-7 minv = 0
+ nfactor = 1.050491 lnfactor = -5.180044E-7 wnfactor = -2.34119E-8
+ pnfactor = 3.269365E-13 eta0 = 0.032 etab = -0.01932
+ dsub = 0.504 cit = -8E-4 cdsc = 0
+ cdscb = 0 cdscd = 0 pclm = -0.821222
+ wpclm = 5.088292E-6 pdiblc1 = 0.21098 pdiblc2 = 2E-4
+ pdiblcb = -0.26831 drout = 0.36075 pscbe1 = 9.3731E8
+ pscbe2 = 1.68E-6 pvag = 1.99 delta = 0.0246
+ fprout = 10.125 pdits = 0 pditsl = 0
+ pditsd = 0 lambda = 0 vtl = 0
+ lc = 5E-9 xn = 3 alpha0 = -7.402317E-6
+ lalpha0 = 9.845692E-11 walpha0 = 6.632109E-11 palpha0 = -3.040897E-16
+ alpha1 = 0 beta0 = 16.919792 lbeta0 = 3.677568E-5
+ wbeta0 = 1.209877E-5 pbeta0 = -4.403409E-11 aigbacc = 1
+ bigbacc = 0 cigbacc = 0 nigbacc = 1
+ aigbinv = 0.35 bigbinv = 0.03 cigbinv = 6E-3
+ eigbinv = 1.1 nigbinv = 3 aigc = 0.43
+ bigc = 0.054 cigc = 0.075 aigsd = 0.43
+ bigsd = 0.054 cigsd = 0.075 dlcig = 0
+ nigc = 1 poxedge = 1 pigcd = 1
+ ntox = 1 toxref = 1.16E-8 agidl = 5.06E-11
+ bgidl = 1.058E9 cgidl = 4E3 egidl = 0.8
+ noia = 2.6E41 noib = 0 noic = 0
+ em = 4.1E7 af = 1 ef = 0.89
+ kf = 0 lintnoi = 0 tnoia = 7.5E6
+ tnoib = 7.2E6 ntnoi = 1 rnoia = 0.794
+ rnoib = 0.38 xpart = 0 cgso = {2.754679E-10/sw_func_tox_hv_ratio}
+ cgdo = {2.754679E-10/sw_func_tox_hv_ratio} cgbo = {0/sw_func_tox_hv_ratio} ckappas = 0.6
+ cf = 0 clc = 1E-7 cle = 0.6
+ dlc = 6.5995E-8 dwc = 0 vfbcv = -1
+ noff = 4 voffcv = -0.4104 acde = 0.4176
+ moin = 15 cgsl = {4.49025E-11/sw_func_tox_hv_ratio} cgdl = {4.49025E-11/sw_func_tox_hv_ratio}
+ ijthsrev = 0.1 ijthsfwd = 0.1 xjbvs = 1
+ bvs = 12.636 jss = 3.75E-4 jsws = 5.84E-11
+ cjs = {8.310E-04*sw_func_nsd_pw_cj} mjs = 0.295 mjsws = 0.037586
+ cjsws = {8.643094E-11*sw_func_nsd_pw_cj} cjswgs = {5.47776E-11*sw_func_nsd_pw_cj} mjswgs = 0.78692
+ pbs = 0.72468 pbsws = 0.29067 pbswgs = 0.54958
+ xrcrg1 = 12 xrcrg2 = 1 rbpb = 50
+ rbpd = 50 rbps = 50 rbdb = 50
+ rbsb = 50 gbmin = 1E-12 tnom = 30
+ ute = -1.33707 lute = 3.018725E-7 kt1 = -0.414271
+ lkt1 = 9.056174E-8 kt1l = 0 kt2 = -0.019151
+ ua1 = 3.0044E-9 ub1 = -3.7525E-18 uc1 = -5.9821E-11
+ at = 3.041925E5 lat = -0.748698 wat = -0.411193
+ pat = 1.017873E-6 prt = 0 njs = 1.0773
+ xtis = 0.76 tpb = 1.344E-3 tpbsw = 9.9005E-4
+ tpbswg = 0 tcj = 6.7434E-4 tcjsw = 2.493E-4
+ tcjswg = 0 tvoff = 0 tvfbsdoff = 0
+ saref = 3E-6 sbref = 3E-6 wlod = 0
+ ku0 = -4.5E-8 kvsat = 0.3 kvth0 = 1.1E-8
+ tku0 = 0 llodku0 = 0 wlodku0 = 1
+ llodvth = 0 wlodvth = 1 lku0 = 0
+ wku0 = 2E-7 pku0 = 0 lkvth0 = 0
+ wkvth0 = 6.5E-7 pkvth0 = 0 stk2 = 0
+ lodk2 = 1 steta0 = 0 lodeta0 = 1

.model nhv_model.31 nmos
+ level = 54 lmin = 2E-6 lmax = 4E-6 wmin = 3E-6
+ wmax = 5E-6 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 1.16E-8
+ toxm = 1.16E-8 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 1E23 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {2.1346E-8+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {7.6507E-8-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = -4.1292E-9 dwb = -1.6944E-9 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = 0.802026 lvth0 = -1.950007E-8
+ wvth0 = -4.463496E-9 pvth0 = 3.37238E-14 k1 = 0.88325
+ k2 = -4.43372E-2 lk2 = 1.400604E-8 wk2 = 1.015567E-8
+ pk2 = 6.898404E-15 k3 = -0.884 k3b = 0.43
+ w0 = 0 lpe0 = 2.5E-8 lpeb = -2.182E-7
+ vbm = -3 dvtp0 = 0 dvtp1 = 0
+ dvt0 = 0 dvt1 = 0.53 dvt2 = -0.19251
+ dvt0w = 0.16 dvt1w = 6.9091E6 dvt2w = -0.036016
+ vfbsdoff = 0 u0 = 4.61562E-2 lu0 = 4.626676E-11
+ wu0 = -1.899176E-8 pu0 = 8.433813E-15 ua = 4.6493E-10
+ lua = -2.902686E-16 wua = -1.810517E-15 pua = 8.512537E-22
+ ub = 1.15786E-18 lub = 2.421204E-25 wub = 1.925137E-24
+ pub = -9.762453E-31 uc = 6.6204E-11 ud = 0
+ up = 0 lp = 1 eu = 1.67
+ vsat = 1.451146E5 lvsat = -6.73472E-2 wvsat = -0.213009
+ pvsat = 3.467171E-7 a0 = 0.177919 la0 = 1.716212E-6
+ wa0 = 1.878507E-6 pa0 = -3.40684E-12 ags = 2.54357E-2
+ lags = 3.437169E-7 wags = 4.764273E-7 pags = -1.143263E-12
+ b0 = 3.2933E-8 b1 = 0 keta = -4.06511E-2
+ lketa = 1.09113E-7 wketa = 3.052273E-8 pketa = -3.226807E-13
+ a1 = 0 a2 = 0.659726 rdsw = 724.62
+ rdswmin = 0 rdw = 0 rdwmin = 0
+ rsw = 0 rswmin = 0 prwb = 0.05626
+ prwg = 0.048 wr = 1 voff = -0.20613
+ voffl = -4.257949E-7 minv = 0 nfactor = 0.956988
+ lnfactor = -1.582998E-7 wnfactor = 5.778238E-8 pnfactor = 1.458326E-14
+ eta0 = 0.032 etab = -0.01932 dsub = 0.504
+ cit = -8E-4 cdsc = 0 cdscb = 0
+ cdscd = 0 pclm = -0.821222 wpclm = 5.088292E-6
+ pdiblc1 = 0.21098 pdiblc2 = 2E-4 pdiblcb = -0.26831
+ drout = 0.36075 pscbe1 = 9.3731E8 pscbe2 = 1.68E-6
+ pvag = 1.99 delta = 0.0246 fprout = 10.125
+ pdits = 0 pditsl = 0 pditsd = 0
+ lambda = 0 vtl = 0 lc = 5E-9
+ xn = 3 alpha0 = 2.162998E-5 lalpha0 = -1.322992E-11
+ walpha0 = -2.44767E-11 palpha0 = 4.520812E-17 alpha1 = 0
+ beta0 = 24.080454 lbeta0 = 9.228711E-6 wbeta0 = -9.925659E-7
+ pbeta0 = 6.328094E-12 aigbacc = 1 bigbacc = 0
+ cigbacc = 0 nigbacc = 1 aigbinv = 0.35
+ bigbinv = 0.03 cigbinv = 6E-3 eigbinv = 1.1
+ nigbinv = 3 aigc = 0.43 bigc = 0.054
+ cigc = 0.075 aigsd = 0.43 bigsd = 0.054
+ cigsd = 0.075 dlcig = 0 nigc = 1
+ poxedge = 1 pigcd = 1 ntox = 1
+ toxref = 1.16E-8 agidl = 5.06E-11 bgidl = 1.058E9
+ cgidl = 4E3 egidl = 0.8 noia = 2.6E41
+ noib = 0 noic = 0 em = 4.1E7
+ af = 1 ef = 0.89 kf = 0
+ lintnoi = 0 tnoia = 7.5E6 tnoib = 7.2E6
+ ntnoi = 1 rnoia = 0.794 rnoib = 0.38
+ xpart = 0 cgso = {2.754679E-10/sw_func_tox_hv_ratio} cgdo = {2.754679E-10/sw_func_tox_hv_ratio}
+ cgbo = {0/sw_func_tox_hv_ratio} ckappas = 0.6 cf = 0
+ clc = 1E-7 cle = 0.6 dlc = 6.5995E-8
+ dwc = 0 vfbcv = -1 noff = 4
+ voffcv = -0.4104 acde = 0.4176 moin = 15
+ cgsl = {4.49025E-11/sw_func_tox_hv_ratio} cgdl = {4.49025E-11/sw_func_tox_hv_ratio} ijthsrev = 0.1
+ ijthsfwd = 0.1 xjbvs = 1 bvs = 12.636
+ jss = 3.75E-4 jsws = 5.84E-11 cjs = {8.310E-04*sw_func_nsd_pw_cj}
+ mjs = 0.295 mjsws = 0.037586 cjsws = {8.643094E-11*sw_func_nsd_pw_cj}
+ cjswgs = {5.47776E-11*sw_func_nsd_pw_cj} mjswgs = 0.78692 pbs = 0.72468
+ pbsws = 0.29067 pbswgs = 0.54958 xrcrg1 = 12
+ xrcrg2 = 1 rbpb = 50 rbpd = 50
+ rbps = 50 rbdb = 50 rbsb = 50
+ gbmin = 1E-12 tnom = 30 ute = -1.22166
+ lute = -1.421066E-7 kt1 = -0.407353 lkt1 = 6.394796E-8
+ kt1l = 0 kt2 = -0.019151 ua1 = 3.0044E-9
+ ub1 = -3.7525E-18 uc1 = -5.9821E-11 at = 1.786379E5
+ lat = -0.265691 wat = -0.214296 pat = 2.604154E-7
+ prt = 0 njs = 1.0773 xtis = 0.76
+ tpb = 1.344E-3 tpbsw = 9.9005E-4 tpbswg = 0
+ tcj = 6.7434E-4 tcjsw = 2.493E-4 tcjswg = 0
+ tvoff = 0 tvfbsdoff = 0 saref = 3E-6
+ sbref = 3E-6 wlod = 0 ku0 = -4.5E-8
+ kvsat = 0.3 kvth0 = 1.1E-8 tku0 = 0
+ llodku0 = 0 wlodku0 = 1 llodvth = 0
+ wlodvth = 1 lku0 = 0 wku0 = 2E-7
+ pku0 = 0 lkvth0 = 0 wkvth0 = 6.5E-7
+ pkvth0 = 0 stk2 = 0 lodk2 = 1
+ steta0 = 0 lodeta0 = 1

.model nhv_model.32 nmos
+ level = 54 lmin = 1E-6 lmax = 2E-6 wmin = 3E-6
+ wmax = 5E-6 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 1.16E-8
+ toxm = 1.16E-8 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 1E23 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {2.1346E-8+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {7.6507E-8-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = -4.1292E-9 dwb = -1.6944E-9 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = 0.80367 lvth0 = -2.253716E-8
+ wvth0 = -4.669437E-8 pvth0 = 1.117236E-13 k1 = 0.88325
+ k2 = -2.61273E-2 lk2 = -1.962743E-8 wk2 = -3.878937E-8
+ pk2 = 9.72992E-14 k3 = -0.884 k3b = 0.43
+ w0 = 0 lpe0 = 2.5E-8 lpeb = -2.182E-7
+ vbm = -3 dvtp0 = 0 dvtp1 = 0
+ dvt0 = 0 dvt1 = 0.53 dvt2 = -0.19251
+ dvt0w = 0.16 dvt1w = 6.9091E6 dvt2w = -0.036016
+ vfbsdoff = 0 u0 = 4.72397E-2 lu0 = -1.955017E-9
+ wu0 = -1.967276E-8 pu0 = 9.69162E-15 ua = 3.088168E-10
+ lua = -1.929873E-18 wua = -1.354809E-15 pua = 9.566973E-24
+ ub = 1.281754E-18 lub = 1.328913E-26 wub = 1.432244E-24
+ pub = -6.587829E-32 uc = 6.6204E-11 ud = 0
+ up = 0 lp = 1 eu = 1.67
+ vsat = 1.099038E5 lvsat = -2.313164E-3 wvsat = -3.14975E-2
+ pvsat = 1.146707E-8 a0 = 1.105428 la0 = 3.114906E-9
+ wa0 = 4.232682E-8 pa0 = -1.544155E-14 ags = 0.216438
+ lags = -9.062513E-9 wags = -1.668848E-7 pags = 4.492567E-14
+ b0 = 3.2933E-8 b1 = 0 keta = 4.30598E-2
+ lketa = -4.549993E-8 wketa = -2.663057E-7 pketa = 2.255572E-13
+ a1 = 0 a2 = 0.659726 rdsw = 724.62
+ rdswmin = 0 rdw = 0 rdwmin = 0
+ rsw = 0 rswmin = 0 prwb = 0.05626
+ prwg = 0.048 wr = 1 voff = -0.20613
+ voffl = -4.257949E-7 minv = 0 nfactor = 0.849477
+ lnfactor = 4.027218E-8 wnfactor = 1.737686E-7 pnfactor = -1.996416E-13
+ eta0 = 0.032 etab = -0.01932 dsub = 0.504
+ cit = -8E-4 cdsc = 0 cdscb = 0
+ cdscd = 0 pclm = -0.821222 wpclm = 5.088292E-6
+ pdiblc1 = 0.21098 pdiblc2 = 2E-4 pdiblcb = -0.26831
+ drout = 0.36075 pscbe1 = 9.3731E8 pscbe2 = 1.68E-6
+ pvag = 1.99 delta = 0.0246 fprout = 10.125
+ pdits = 0 pditsl = 0 pditsd = 0
+ lambda = 0 vtl = 0 lc = 5E-9
+ xn = 3 alpha0 = 1.990241E-5 lalpha0 = -1.003913E-11
+ walpha0 = -2.694501E-11 palpha0 = 4.976707E-17 alpha1 = 0
+ beta0 = 34.215681 lbeta0 = -9.490911E-6 wbeta0 = -2.303999E-5
+ pbeta0 = 4.704937E-11 aigbacc = 1 bigbacc = 0
+ cigbacc = 0 nigbacc = 1 aigbinv = 0.35
+ bigbinv = 0.03 cigbinv = 6E-3 eigbinv = 1.1
+ nigbinv = 3 aigc = 0.43 bigc = 0.054
+ cigc = 0.075 aigsd = 0.43 bigsd = 0.054
+ cigsd = 0.075 dlcig = 0 nigc = 1
+ poxedge = 1 pigcd = 1 ntox = 1
+ toxref = 1.16E-8 agidl = 5.06E-11 bgidl = 1.058E9
+ cgidl = 4E3 egidl = 0.8 noia = 2.6E41
+ noib = 0 noic = 0 em = 4.1E7
+ af = 1 ef = 0.89 kf = 0
+ lintnoi = 0 tnoia = 7.5E6 tnoib = 7.2E6
+ ntnoi = 1 rnoia = 0.794 rnoib = 0.38
+ xpart = 0 cgso = {2.754679E-10/sw_func_tox_hv_ratio} cgdo = {2.754679E-10/sw_func_tox_hv_ratio}
+ cgbo = {0/sw_func_tox_hv_ratio} ckappas = 0.6 cf = 0
+ clc = 1E-7 cle = 0.6 dlc = 6.5995E-8
+ dwc = 0 vfbcv = -1 noff = 4
+ voffcv = -0.4104 acde = 0.4176 moin = 15
+ cgsl = {4.49025E-11/sw_func_tox_hv_ratio} cgdl = {4.49025E-11/sw_func_tox_hv_ratio} ijthsrev = 0.1
+ ijthsfwd = 0.1 xjbvs = 1 bvs = 12.636
+ jss = 3.75E-4 jsws = 5.84E-11 cjs = {8.310E-04*sw_func_nsd_pw_cj}
+ mjs = 0.295 mjsws = 0.037586 cjsws = {8.643094E-11*sw_func_nsd_pw_cj}
+ cjswgs = {5.47776E-11*sw_func_nsd_pw_cj} mjswgs = 0.78692 pbs = 0.72468
+ pbsws = 0.29067 pbswgs = 0.54958 xrcrg1 = 12
+ xrcrg2 = 1 rbpb = 50 rbpd = 50
+ rbps = 50 rbdb = 50 rbsb = 50
+ gbmin = 1E-12 tnom = 30 ute = -1.2986
+ kt1 = -0.37273 kt1l = 0 kt2 = -0.019151
+ ua1 = 3.0044E-9 ub1 = -3.37678E-18 lub1 = -6.939492E-25
+ wub1 = -1.862559E-24 pub1 = 3.44012E-30 uc1 = -5.9821E-11
+ at = 5.232013E4 lat = -3.23843E-2 wat = -0.160221
+ pat = 1.605389E-7 prt = 0 njs = 1.0773
+ xtis = 0.76 tpb = 1.344E-3 tpbsw = 9.9005E-4
+ tpbswg = 0 tcj = 6.7434E-4 tcjsw = 2.493E-4
+ tcjswg = 0 tvoff = 0 tvfbsdoff = 0
+ saref = 3E-6 sbref = 3E-6 wlod = 0
+ ku0 = -4.5E-8 kvsat = 0.3 kvth0 = 1.1E-8
+ tku0 = 0 llodku0 = 0 wlodku0 = 1
+ llodvth = 0 wlodvth = 1 lku0 = 0
+ wku0 = 2E-7 pku0 = 0 lkvth0 = 0
+ wkvth0 = 6.5E-7 pkvth0 = 0 stk2 = 0
+ lodk2 = 1 steta0 = 0 lodeta0 = 1

.model nhv_model.33 nmos
+ level = 54 lmin = 8E-7 lmax = 1E-6 wmin = 3E-6
+ wmax = 5E-6 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 1.16E-8
+ toxm = 1.16E-8 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 1E23 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {2.1346E-8+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {7.6507E-8-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = -4.1292E-9 dwb = -1.6944E-9 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = 0.686904 lvth0 = 7.63621E-8
+ wvth0 = 3.518363E-7 pvth0 = -2.258262E-13 k1 = 0.88325
+ k2 = -0.067057 lk2 = 1.503948E-8 wk2 = 1.28599E-7
+ pk2 = -4.447636E-14 k3 = -0.884 k3b = 0.43
+ w0 = 0 lpe0 = 2.5E-8 lpeb = -2.182E-7
+ vbm = -3 dvtp0 = 0 dvtp1 = 0
+ dvt0 = 0 dvt1 = 0.53 dvt2 = -0.19251
+ dvt0w = 0.16 dvt1w = 6.9091E6 dvt2w = -0.036016
+ vfbsdoff = 0 u0 = 3.696766E-3 lu0 = 3.492527E-8
+ wu0 = 1.137136E-7 pu0 = -1.032848E-13 ua = 1.78684E-9
+ lua = -1.253795E-15 wua = -5.721223E-15 pua = 3.707859E-21
+ ub = -9.524417E-18 lub = 9.165965E-24 wub = 3.335804E-23
+ pub = -2.710658E-29 uc = 6.6204E-11 ud = 0
+ up = 0 lp = 1 eu = 1.67
+ vsat = 8.937935E4 lvsat = 1.50707E-2 wvsat = 3.46616E-2
+ pvsat = -4.456875E-8 a0 = 1.043089 la0 = 5.591534E-8
+ wa0 = 2.193278E-7 pa0 = -1.653589E-13 ags = 0.386342
+ lags = -1.529687E-7 wags = -6.479434E-7 pags = 4.523755E-13
+ b0 = 3.2933E-8 b1 = 0 keta = -0.01066
+ a1 = 0 a2 = 0.659726 rdsw = 724.62
+ rdswmin = 0 rdw = 0 rdwmin = 0
+ rsw = 0 rswmin = 0 prwb = 0.05626
+ prwg = 0.048 wr = 1 voff = -0.20613
+ voffl = -4.257949E-7 minv = 0 nfactor = 1.558131
+ lnfactor = -5.59948E-7 wnfactor = -2.017035E-6 pnfactor = 1.655939E-12
+ eta0 = 0.032 etab = -0.01932 dsub = 0.504
+ cit = -8E-4 cdsc = 0 cdscb = 0
+ cdscd = 0 pclm = -9.477749 lpclm = 7.331957E-6
+ wpclm = 3.068831E-5 ppclm = -2.168285E-11 pdiblc1 = 0.21098
+ pdiblc2 = 2E-4 pdiblcb = -0.26831 drout = 0.36075
+ pscbe1 = 9.3731E8 pscbe2 = 1.68E-6 pvag = 1.99
+ delta = 0.0246 fprout = 10.125 pdits = 0
+ pditsl = 0 pditsd = 0 lambda = 0
+ vtl = 0 lc = 5E-9 xn = 3
+ alpha0 = 8.049642E-6 walpha0 = 3.181282E-11 alpha1 = 0
+ beta0 = -36.260898 lbeta0 = 5.020176E-5 wbeta0 = 2.07792E-4
+ pbeta0 = -1.484621E-10 aigbacc = 1 bigbacc = 0
+ cigbacc = 0 nigbacc = 1 aigbinv = 0.35
+ bigbinv = 0.03 cigbinv = 6E-3 eigbinv = 1.1
+ nigbinv = 3 aigc = 0.43 bigc = 0.054
+ cigc = 0.075 aigsd = 0.43 bigsd = 0.054
+ cigsd = 0.075 dlcig = 0 nigc = 1
+ poxedge = 1 pigcd = 1 ntox = 1
+ toxref = 1.16E-8 agidl = 5.06E-11 bgidl = 1.058E9
+ cgidl = 4E3 egidl = 0.8 noia = 2.6E41
+ noib = 0 noic = 0 em = 4.1E7
+ af = 1 ef = 0.89 kf = 0
+ lintnoi = 0 tnoia = 7.5E6 tnoib = 7.2E6
+ ntnoi = 1 rnoia = 0.794 rnoib = 0.38
+ xpart = 0 cgso = {2.754679E-10/sw_func_tox_hv_ratio} cgdo = {2.754679E-10/sw_func_tox_hv_ratio}
+ cgbo = {0/sw_func_tox_hv_ratio} ckappas = 0.6 cf = 0
+ clc = 1E-7 cle = 0.6 dlc = 6.5995E-8
+ dwc = 0 vfbcv = -1 noff = 4
+ voffcv = -0.4104 acde = 0.4176 moin = 15
+ cgsl = {4.49025E-11/sw_func_tox_hv_ratio} cgdl = {4.49025E-11/sw_func_tox_hv_ratio} ijthsrev = 0.1
+ ijthsfwd = 0.1 xjbvs = 1 bvs = 12.636
+ jss = 3.75E-4 jsws = 5.84E-11 cjs = {8.310E-04*sw_func_nsd_pw_cj}
+ mjs = 0.295 mjsws = 0.037586 cjsws = {8.643094E-11*sw_func_nsd_pw_cj}
+ cjswgs = {5.47776E-11*sw_func_nsd_pw_cj} mjswgs = 0.78692 pbs = 0.72468
+ pbsws = 0.29067 pbswgs = 0.54958 xrcrg1 = 12
+ xrcrg2 = 1 rbpb = 50 rbpd = 50
+ rbps = 50 rbdb = 50 rbsb = 50
+ gbmin = 1E-12 tnom = 30 ute = -1.2986
+ kt1 = -0.549132 lkt1 = 1.4941E-7 wkt1 = 5.21675E-7
+ pkt1 = -4.418514E-13 kt1l = 0 kt2 = -0.019151
+ ua1 = 3.0044E-9 ub1 = -5.799751E-18 lub1 = 1.358273E-24
+ wub1 = 6.941543E-24 pub1 = -4.016831E-30 uc1 = -5.9821E-11
+ at = -2.232555E5 lat = 0.201024 wat = 0.731211
+ pat = -5.94491E-7 prt = 0 njs = 1.0773
+ xtis = 0.76 tpb = 1.344E-3 tpbsw = 9.9005E-4
+ tpbswg = 0 tcj = 6.7434E-4 tcjsw = 2.493E-4
+ tcjswg = 0 tvoff = 0 tvfbsdoff = 0
+ saref = 2.81E-6 sbref = 2.81E-6 wlod = 0
+ ku0 = -4.5E-8 kvsat = 0.3 kvth0 = 1.1E-8
+ tku0 = 0 llodku0 = 0 wlodku0 = 1
+ llodvth = 0 wlodvth = 1 lku0 = 0
+ wku0 = 2E-7 pku0 = 0 lkvth0 = 0
+ wkvth0 = 6.5E-7 pkvth0 = 0 stk2 = 0
+ lodk2 = 1 steta0 = 0 lodeta0 = 1

.model nhv_model.34 nmos
+ level = 54 lmin = 6E-7 lmax = 8E-7 wmin = 3E-6
+ wmax = 5E-6 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 1.16E-8
+ toxm = 1.16E-8 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 1E23 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {2.1346E-8+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {7.6507E-8-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = -4.1292E-9 dwb = -1.6944E-9 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = 0.862615 lvth0 = -3.732031E-8
+ wvth0 = -2.831613E-7 pvth0 = 1.850083E-13 k1 = 0.88325
+ k2 = -4.74629E-2 lk2 = 2.362372E-9 wk2 = 7.795588E-8
+ pk2 = -1.171101E-14 k3 = -0.884 k3b = 0.43
+ w0 = 0 lpe0 = 2.5E-8 lpeb = -2.182E-7
+ vbm = -3 dvtp0 = 0 dvtp1 = 0
+ dvt0 = 0 dvt1 = 0.53 dvt2 = -0.19251
+ dvt0w = 0.16 dvt1w = 6.9091E6 dvt2w = -0.036016
+ vfbsdoff = 0 u0 = 6.78868E-2 lu0 = -6.604765E-9
+ wu0 = -9.653302E-8 pu0 = 3.274185E-14 ua = -1.475823E-10
+ lua = -2.250764E-18 wua = -7.496617E-18 pua = 1.115773E-23
+ ub = 6.711957E-18 lub = -1.338742E-24 wub = -1.879631E-23
+ pub = 6.636555E-30 uc = 6.6204E-11 ud = 0
+ up = 0 lp = 1 eu = 1.67
+ vsat = 1.158717E5 lvsat = -2.069454E-3 wvsat = -5.00817E-2
+ pvsat = 1.025892E-8 a0 = 1.145859 la0 = -1.057519E-8
+ wa0 = -1.172844E-7 pa0 = 5.242448E-14 ags = 0.126799
+ lags = 1.495207E-8 wags = 1.658263E-7 pags = -7.412202E-14
+ b0 = 3.2933E-8 b1 = 0 keta = -0.01066
+ a1 = 0 a2 = 0.659726 rdsw = 724.62
+ rdswmin = 0 rdw = 0 rdwmin = 0
+ rsw = 0 rswmin = 0 prwb = 0.05626
+ prwg = 0.048 wr = 1 voff = -0.20613
+ voffl = -4.257949E-7 minv = 0 nfactor = 0.566718
+ lnfactor = 8.14825E-8 wnfactor = 1.166762E-6 pnfactor = -4.039338E-13
+ eta0 = 0.032 etab = -0.01932 dsub = 0.504
+ cit = -8E-4 cdsc = 0 cdscb = 0
+ cdscd = 0 pclm = 3.128491 lpclm = -8.241042E-7
+ wpclm = -9.139746E-6 ppclm = 4.085339E-12 pdiblc1 = 0.21098
+ pdiblc2 = 2E-4 pdiblcb = -0.26831 drout = 0.36075
+ pscbe1 = 9.3731E8 pscbe2 = 1.68E-6 pvag = 1.99
+ delta = 0.0246 fprout = 10.125 pdits = 0
+ pditsl = 0 pditsd = 0 lambda = 0
+ vtl = 0 lc = 5E-9 xn = 3
+ alpha0 = 6.136227E-6 lalpha0 = 1.237952E-12 walpha0 = 4.129821E-11
+ palpha0 = -6.136911E-18 alpha1 = 0 beta0 = 51.104343
+ lbeta0 = -6.322323E-6 wbeta0 = -7.011786E-5 pbeta0 = 3.13417E-11
+ aigbacc = 1 bigbacc = 0 cigbacc = 0
+ nigbacc = 1 aigbinv = 0.35 bigbinv = 0.03
+ cigbinv = 6E-3 eigbinv = 1.1 nigbinv = 3
+ aigc = 0.43 bigc = 0.054 cigc = 0.075
+ aigsd = 0.43 bigsd = 0.054 cigsd = 0.075
+ dlcig = 0 nigc = 1 poxedge = 1
+ pigcd = 1 ntox = 1 toxref = 1.16E-8
+ agidl = 5.06E-11 bgidl = 1.058E9 cgidl = 4E3
+ egidl = 0.8 noia = 2.6E41 noib = 0
+ noic = 0 em = 4.1E7 af = 1
+ ef = 0.89 kf = 0 lintnoi = 0
+ tnoia = 7.5E6 tnoib = 7.2E6 ntnoi = 1
+ rnoia = 0.794 rnoib = 0.38 xpart = 0
+ cgso = {2.754679E-10/sw_func_tox_hv_ratio} cgdo = {2.754679E-10/sw_func_tox_hv_ratio} cgbo = {0/sw_func_tox_hv_ratio}
+ ckappas = 0.6 cf = 0 clc = 1E-7
+ cle = 0.6 dlc = 6.5995E-8 dwc = 0
+ vfbcv = -1 noff = 4 voffcv = -0.4104
+ acde = 0.4176 moin = 15 cgsl = {4.49025E-11/sw_func_tox_hv_ratio}
+ cgdl = {4.49025E-11/sw_func_tox_hv_ratio} ijthsrev = 0.1 ijthsfwd = 0.1
+ xjbvs = 1 bvs = 12.636 jss = 3.75E-4
+ jsws = 5.84E-11 cjs = {8.310E-04*sw_func_nsd_pw_cj} mjs = 0.295
+ mjsws = 0.037586 cjsws = {8.643094E-11*sw_func_nsd_pw_cj} cjswgs = {5.47776E-11*sw_func_nsd_pw_cj}
+ mjswgs = 0.78692 pbs = 0.72468 pbsws = 0.29067
+ pbswgs = 0.54958 xrcrg1 = 12 xrcrg2 = 1
+ rbpb = 50 rbpd = 50 rbps = 50
+ rbdb = 50 rbsb = 50 gbmin = 1E-12
+ tnom = 30 ute = -1.2986 kt1 = -0.31159
+ lkt1 = -4.276174E-9 wkt1 = -1.940279E-7 pkt1 = 2.119831E-14
+ kt1l = 0 kt2 = -0.019151 ua1 = -2.76164E-10
+ lua1 = 2.122479E-15 wua1 = 1.626277E-14 pua1 = -1.052178E-20
+ ub1 = 2.709077E-18 lub1 = -4.14682E-24 wub1 = -3.104057E-23
+ pub1 = 2.055706E-29 uc1 = -5.9821E-11 at = 1.350411E5
+ lat = -3.07885E-2 wat = -0.423558 pat = 1.526278E-7
+ prt = 0 njs = 1.0773 xtis = 0.76
+ tpb = 1.344E-3 tpbsw = 9.9005E-4 tpbswg = 0
+ tcj = 6.7434E-4 tcjsw = 2.493E-4 tcjswg = 0
+ tvoff = 0 tvfbsdoff = 0 saref = 2.81E-6
+ sbref = 2.81E-6 wlod = 0 ku0 = -4.5E-8
+ kvsat = 0.3 kvth0 = 1.1E-8 tku0 = 0
+ llodku0 = 0 wlodku0 = 1 llodvth = 0
+ wlodvth = 1 lku0 = 0 wku0 = 2E-7
+ pku0 = 0 lkvth0 = 0 wkvth0 = 6.5E-7
+ pkvth0 = 0 stk2 = 0 lodk2 = 1
+ steta0 = 0 lodeta0 = 1

.model nhv_model.35 nmos
+ level = 54 lmin = 5E-7 lmax = 6E-7 wmin = 3E-6
+ wmax = 5E-6 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 1.16E-8
+ toxm = 1.16E-8 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 1E23 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {2.1346E-8+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {7.6507E-8-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = -4.1292E-9 dwb = -1.6944E-9 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = 0.714588 lvth0 = 2.88459E-8
+ wvth0 = 4.506565E-7 pvth0 = -1.42998E-13 k1 = 0.88325
+ k2 = -7.11957E-2 lk2 = 1.297056E-8 wk2 = 1.956062E-7
+ pk2 = -6.429907E-14 k3 = -0.884 k3b = 0.43
+ w0 = 0 lpe0 = 2.5E-8 lpeb = -2.182E-7
+ vbm = -3 dvtp0 = 0 dvtp1 = 0
+ dvt0 = 0 dvt1 = 0.53 dvt2 = -0.19251
+ dvt0w = 0.16 dvt1w = 6.9091E6 dvt2w = -0.036016
+ vfbsdoff = 0 u0 = 6.24223E-2 lu0 = -4.162221E-9
+ wu0 = -6.944394E-8 pu0 = 2.063341E-14 ua = -1.531272E-10
+ lua = 2.277308E-19 wua = 1.999119E-17 pua = -1.128931E-24
+ ub = 5.94565E-18 lub = -9.962131E-25 wub = -1.499749E-23
+ pub = 4.938535E-30 uc = 6.6204E-11 ud = 0
+ up = 0 lp = 1 eu = 1.67
+ vsat = 1.404424E5 lvsat = -1.30522E-2 wvsat = -0.171886
+ pvsat = 6.47038E-8 a0 = 1.1222 ags = 0.16025
+ b0 = 3.2933E-8 b1 = 0 keta = -0.01066
+ a1 = 0 a2 = 0.659726 rdsw = 724.62
+ rdswmin = 0 rdw = 0 rdwmin = 0
+ rsw = 0 rswmin = 0 prwb = 0.05626
+ prwg = 0.048 wr = 1 voff = -0.20613
+ voffl = -4.257949E-7 minv = 0 nfactor = 0.911604
+ lnfactor = -7.267661E-8 wnfactor = -5.429427E-7 pnfactor = 3.602804E-13
+ eta0 = 0.032 etab = -0.01932 dsub = 0.504
+ cit = -8E-4 cdsc = 0 cdscb = 0
+ cdscd = 0 pclm = 1.2848 pdiblc1 = 0.21098
+ pdiblc2 = 2E-4 pdiblcb = -0.26831 drout = 0.36075
+ pscbe1 = 9.3731E8 pscbe2 = 1.68E-6 pvag = 1.99
+ delta = 0.0246 fprout = 10.125 pdits = 0
+ pditsl = 0 pditsd = 0 lambda = 0
+ vtl = 0 lc = 5E-9 xn = 3
+ alpha0 = -1.039086E-5 lalpha0 = 8.625331E-12 walpha0 = 1.232281E-10
+ palpha0 = -4.275842E-17 alpha1 = 0 beta0 = 36.96
+ aigbacc = 1 bigbacc = 0 cigbacc = 0
+ nigbacc = 1 aigbinv = 0.35 bigbinv = 0.03
+ cigbinv = 6E-3 eigbinv = 1.1 nigbinv = 3
+ aigc = 0.43 bigc = 0.054 cigc = 0.075
+ aigsd = 0.43 bigsd = 0.054 cigsd = 0.075
+ dlcig = 0 nigc = 1 poxedge = 1
+ pigcd = 1 ntox = 1 toxref = 1.16E-8
+ agidl = 5.06E-11 bgidl = 1.058E9 cgidl = 4E3
+ egidl = 0.8 noia = 2.6E41 noib = 0
+ noic = 0 em = 4.1E7 af = 1
+ ef = 0.89 kf = 0 lintnoi = 0
+ tnoia = 7.5E6 tnoib = 7.2E6 ntnoi = 1
+ rnoia = 0.794 rnoib = 0.38 xpart = 0
+ cgso = {2.754679E-10/sw_func_tox_hv_ratio} cgdo = {2.754679E-10/sw_func_tox_hv_ratio} cgbo = {0/sw_func_tox_hv_ratio}
+ ckappas = 0.6 cf = 0 clc = 1E-7
+ cle = 0.6 dlc = 6.5995E-8 dwc = 0
+ vfbcv = -1 noff = 4 voffcv = -0.4104
+ acde = 0.4176 moin = 15 cgsl = {4.49025E-11/sw_func_tox_hv_ratio}
+ cgdl = {4.49025E-11/sw_func_tox_hv_ratio} ijthsrev = 0.1 ijthsfwd = 0.1
+ xjbvs = 1 bvs = 12.636 jss = 3.75E-4
+ jsws = 5.84E-11 cjs = {8.310E-04*sw_func_nsd_pw_cj} mjs = 0.295
+ mjsws = 0.037586 cjsws = {8.643094E-11*sw_func_nsd_pw_cj} cjswgs = {5.47776E-11*sw_func_nsd_pw_cj}
+ mjswgs = 0.78692 pbs = 0.72468 pbsws = 0.29067
+ pbswgs = 0.54958 xrcrg1 = 12 xrcrg2 = 1
+ rbpb = 50 rbpd = 50 rbps = 50
+ rbdb = 50 rbsb = 50 gbmin = 1E-12
+ tnom = 30 ute = -1.2991 kt1 = -0.218542
+ lkt1 = -4.586722E-8 wkt1 = -6.552943E-7 pkt1 = 2.273779E-13
+ kt1l = 0 kt2 = -0.019151 ua1 = 9.565528E-9
+ lua1 = -2.27662E-15 wua1 = -3.252553E-14 pua1 = 1.12859E-20
+ ub1 = -1.703232E-17 lub1 = 4.67731E-24 wub1 = 6.682363E-23
+ pub1 = -2.318687E-29 uc1 = -5.9821E-11 at = 1.23625E5
+ lat = -2.56856E-2 wat = -0.366965 pat = 1.273316E-7
+ prt = 0 njs = 1.0773 xtis = 0.76
+ tpb = 1.344E-3 tpbsw = 9.9005E-4 tpbswg = 0
+ tcj = 6.7434E-4 tcjsw = 2.493E-4 tcjswg = 0
+ tvoff = 0 tvfbsdoff = 0 saref = 2.02E-6
+ sbref = 2.01E-6 wlod = 0 ku0 = -4.5E-8
+ kvsat = 0.3 kvth0 = 1.1E-8 tku0 = 0
+ llodku0 = 0 wlodku0 = 1 llodvth = 0
+ wlodvth = 1 lku0 = 0 wku0 = 2E-7
+ pku0 = 0 lkvth0 = 0 wkvth0 = 6.5E-7
+ pkvth0 = 0 stk2 = 0 lodk2 = 1
+ steta0 = 0 lodeta0 = 1

.model nhv_model.36 nmos
+ level = 54 lmin = 8E-6 lmax = 2.02E-5 wmin = 1E-6
+ wmax = 3E-6 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 1.16E-8
+ toxm = 1.16E-8 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 1E23 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {2.1346E-8+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {7.6507E-8-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = -4.1292E-9 dwb = -1.6944E-9 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = 0.791079 wvth0 = 1.298746E-8
+ k1 = 0.88325 k2 = -3.90488E-2 wk2 = 2.004387E-9
+ k3 = -0.884 k3b = 0.43 w0 = 0
+ lpe0 = 2.5E-8 lpeb = -2.182E-7 vbm = -3
+ dvtp0 = 0 dvtp1 = 0 dvt0 = 0
+ dvt1 = 0.53 dvt2 = -0.19251 dvt0w = 0.16
+ dvt1w = 6.9091E6 dvt2w = -0.036016 vfbsdoff = 0
+ u0 = 4.12898E-2 wu0 = -2.61891E-9 ua = -1.477251E-10
+ wua = -7.258824E-19 ub = 1.771673E-18 wub = 1.072828E-26
+ uc = 7.269359E-11 wuc = -1.919172E-17 ud = 0
+ up = 0 lp = 1 eu = 1.67
+ vsat = 6.180912E4 wvsat = 4.79524E-2 a0 = 0.885783
+ wa0 = 2.259057E-7 ags = 0.166008 wags = -6.743855E-9
+ b0 = 3.2933E-8 b1 = 0 keta = -3.43947E-2
+ wketa = 1.202066E-8 a1 = 0 a2 = 0.659726
+ rdsw = 724.62 rdswmin = 0 rdw = 0
+ rdwmin = 0 rsw = 0 rswmin = 0
+ prwb = 0.05626 prwg = 0.048 wr = 1
+ voff = -0.20613 voffl = -4.257949E-7 minv = 0
+ nfactor = 0.946059 wnfactor = 1.318705E-7 eta0 = 0.032
+ etab = -0.01932 dsub = 0.504 cit = -8E-4
+ cdsc = 0 cdscb = 0 cdscd = 0
+ pclm = 0.837882 wpclm = 1.818103E-7 pdiblc1 = 0.21098
+ pdiblc2 = 2E-4 pdiblcb = -0.26831 drout = 0.36075
+ pscbe1 = 9.3731E8 pscbe2 = 1.68E-6 pvag = 1.99
+ delta = 0.0246 fprout = 10.125 pdits = 0
+ pditsl = 0 pditsd = 0 lambda = 0
+ vtl = 0 lc = 5E-9 xn = 3
+ alpha0 = 6.641964E-6 walpha0 = 2.314104E-11 alpha1 = 0
+ beta0 = 22.284581 wbeta0 = 4.481559E-6 aigbacc = 1
+ bigbacc = 0 cigbacc = 0 nigbacc = 1
+ aigbinv = 0.35 bigbinv = 0.03 cigbinv = 6E-3
+ eigbinv = 1.1 nigbinv = 3 aigc = 0.43
+ bigc = 0.054 cigc = 0.075 aigsd = 0.43
+ bigsd = 0.054 cigsd = 0.075 dlcig = 0
+ nigc = 1 poxedge = 1 pigcd = 1
+ ntox = 1 toxref = 1.16E-8 agidl = 5.06E-11
+ bgidl = 1.058E9 cgidl = 4E3 egidl = 0.8
+ noia = 2.6E41 noib = 0 noic = 0
+ em = 4.1E7 af = 1 ef = 0.89
+ kf = 0 lintnoi = 0 tnoia = 7.5E6
+ tnoib = 7.2E6 ntnoi = 1 rnoia = 0.794
+ rnoib = 0.38 xpart = 0 cgso = {2.754679E-10/sw_func_tox_hv_ratio}
+ cgdo = {2.754679E-10/sw_func_tox_hv_ratio} cgbo = {0/sw_func_tox_hv_ratio} ckappas = 0.6
+ cf = 0 clc = 1E-7 cle = 0.6
+ dlc = 6.5995E-8 dwc = 0 vfbcv = -1
+ noff = 4 voffcv = -0.4104 acde = 0.4176
+ moin = 15 cgsl = {4.49025E-11/sw_func_tox_hv_ratio} cgdl = {4.49025E-11/sw_func_tox_hv_ratio}
+ ijthsrev = 0.1 ijthsfwd = 0.1 xjbvs = 1
+ bvs = 12.636 jss = 3.75E-4 jsws = 5.84E-11
+ cjs = {8.310E-04*sw_func_nsd_pw_cj} mjs = 0.295 mjsws = 0.037586
+ cjsws = {8.643094E-11*sw_func_nsd_pw_cj} cjswgs = {5.47776E-11*sw_func_nsd_pw_cj} mjswgs = 0.78692
+ pbs = 0.72468 pbsws = 0.29067 pbswgs = 0.54958
+ xrcrg1 = 12 xrcrg2 = 1 rbpb = 50
+ rbpd = 50 rbps = 50 rbdb = 50
+ rbsb = 50 gbmin = 1E-12 tnom = 30
+ ute = -1.360777 wute = 1.83877E-7 kt1 = -0.407517
+ wkt1 = 1.415527E-8 kt1l = 0 kt2 = -0.019151
+ ua1 = 3.0044E-9 ub1 = -3.7525E-18 uc1 = -5.9821E-11
+ at = 9.617699E4 wat = 5.15252E-2 prt = 0
+ njs = 1.0773 xtis = 0.76 tpb = 1.344E-3
+ tpbsw = 9.9005E-4 tpbswg = 0 tcj = 6.7434E-4
+ tcjsw = 2.493E-4 tcjswg = 0 tvoff = 0
+ tvfbsdoff = 0 saref = 3E-6 sbref = 3E-6
+ wlod = 0 ku0 = -4.5E-8 kvsat = 0.3
+ kvth0 = 1.1E-8 tku0 = 0 llodku0 = 0
+ wlodku0 = 1 llodvth = 0 wlodvth = 1
+ lku0 = 0 wku0 = 2E-7 pku0 = 0
+ lkvth0 = 0 wkvth0 = 6.5E-7 pkvth0 = 0
+ stk2 = 0 lodk2 = 1 steta0 = 0
+ lodeta0 = 1

.model nhv_model.37 nmos
+ level = 54 lmin = 4E-6 lmax = 8E-6 wmin = 1E-6
+ wmax = 3E-6 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 1.16E-8
+ toxm = 1.16E-8 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 1E23 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {2.1346E-8+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {7.6507E-8-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = -4.1292E-9 dwb = -1.6944E-9 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = 0.787659 lvth0 = 2.683699E-8
+ wvth0 = 1.473683E-8 pvth0 = -1.372729E-14 k1 = 0.88325
+ k2 = -4.05734E-2 lk2 = 1.196348E-8 wk2 = 1.635317E-9
+ pk2 = 2.896085E-15 k3 = -0.884 k3b = 0.43
+ w0 = 0 lpe0 = 2.5E-8 lpeb = -2.182E-7
+ vbm = -3 dvtp0 = 0 dvtp1 = 0
+ dvt0 = 0 dvt1 = 0.53 dvt2 = -0.19251
+ dvt0w = 0.16 dvt1w = 6.9091E6 dvt2w = -0.036016
+ vfbsdoff = 0 u0 = 4.12786E-2 lu0 = 8.817174E-11
+ wu0 = -2.8226E-9 pu0 = 1.598359E-15 ua = -1.473051E-10
+ lua = -3.296039E-18 wua = -2.119662E-18 pua = 1.093697E-23
+ ub = 1.775426E-18 lub = -2.945131E-26 wub = -3.069574E-26
+ pub = 3.250537E-31 uc = 7.269359E-11 wuc = -1.919172E-17
+ ud = 0 up = 0 lp = 1
+ eu = 1.67 vsat = 5.038689E4 lvsat = 0.08963
+ wvsat = 0.058887 pvsat = -8.580359E-8 a0 = 0.887824
+ la0 = -1.601928E-8 wa0 = 2.266465E-7 pa0 = -5.81268E-15
+ ags = 0.154387 lags = 9.11958E-8 wags = -5.552377E-9
+ pags = -9.349514E-15 b0 = 3.2933E-8 b1 = 0
+ keta = -3.43947E-2 wketa = 1.202066E-8 a1 = 0
+ a2 = 0.659726 rdsw = 724.62 rdswmin = 0
+ rdw = 0 rdwmin = 0 rsw = 0
+ rswmin = 0 prwb = 0.05626 prwg = 0.048
+ wr = 1 voff = -0.20613 voffl = -4.257949E-7
+ minv = 0 nfactor = 0.991713 lnfactor = -3.582527E-7
+ wnfactor = 1.504125E-7 pnfactor = -1.454986E-13 eta0 = 0.032
+ etab = -0.01932 dsub = 0.504 cit = -8E-4
+ cdsc = 0 cdscb = 0 cdscd = 0
+ pclm = 0.837882 wpclm = 1.818103E-7 pdiblc1 = 0.21098
+ pdiblc2 = 2E-4 pdiblcb = -0.26831 drout = 0.36075
+ pscbe1 = 9.3731E8 pscbe2 = 1.68E-6 pvag = 1.99
+ delta = 0.0246 fprout = 10.125 pdits = 0
+ pditsl = 0 pditsd = 0 lambda = 0
+ vtl = 0 lc = 5E-9 xn = 3
+ alpha0 = 3.269781E-6 lalpha0 = 2.646147E-11 walpha0 = 3.476041E-11
+ palpha0 = -9.117699E-17 alpha1 = 0 beta0 = 18.677946
+ lbeta0 = 2.830122E-5 wbeta0 = 6.899368E-6 pbeta0 = -1.897251E-11
+ aigbacc = 1 bigbacc = 0 cigbacc = 0
+ nigbacc = 1 aigbinv = 0.35 bigbinv = 0.03
+ cigbinv = 6E-3 eigbinv = 1.1 nigbinv = 3
+ aigc = 0.43 bigc = 0.054 cigc = 0.075
+ aigsd = 0.43 bigsd = 0.054 cigsd = 0.075
+ dlcig = 0 nigc = 1 poxedge = 1
+ pigcd = 1 ntox = 1 toxref = 1.16E-8
+ agidl = 5.06E-11 bgidl = 1.058E9 cgidl = 4E3
+ egidl = 0.8 noia = 2.6E41 noib = 0
+ noic = 0 em = 4.1E7 af = 1
+ ef = 0.89 kf = 0 lintnoi = 0
+ tnoia = 7.5E6 tnoib = 7.2E6 ntnoi = 1
+ rnoia = 0.794 rnoib = 0.38 xpart = 0
+ cgso = {2.754679E-10/sw_func_tox_hv_ratio} cgdo = {2.754679E-10/sw_func_tox_hv_ratio} cgbo = {0/sw_func_tox_hv_ratio}
+ ckappas = 0.6 cf = 0 clc = 1E-7
+ cle = 0.6 dlc = 6.5995E-8 dwc = 0
+ vfbcv = -1 noff = 4 voffcv = -0.4104
+ acde = 0.4176 moin = 15 cgsl = {4.49025E-11/sw_func_tox_hv_ratio}
+ cgdl = {4.49025E-11/sw_func_tox_hv_ratio} ijthsrev = 0.1 ijthsfwd = 0.1
+ xjbvs = 1 bvs = 12.636 jss = 3.75E-4
+ jsws = 5.84E-11 cjs = {8.310E-04*sw_func_nsd_pw_cj} mjs = 0.295
+ mjsws = 0.037586 cjsws = {8.643094E-11*sw_func_nsd_pw_cj} cjswgs = {5.47776E-11*sw_func_nsd_pw_cj}
+ mjswgs = 0.78692 pbs = 0.72468 pbsws = 0.29067
+ pbswgs = 0.54958 xrcrg1 = 12 xrcrg2 = 1
+ rbpb = 50 rbpd = 50 rbps = 50
+ rbdb = 50 rbsb = 50 gbmin = 1E-12
+ tnom = 30 ute = -1.417661 lute = 4.463649E-7
+ wute = 2.383321E-7 pute = -4.273087E-13 kt1 = -0.423661
+ lkt1 = 1.266849E-7 wkt1 = 2.776906E-8 pkt1 = -1.068272E-13
+ kt1l = 0 kt2 = -0.019151 ua1 = 3.0044E-9
+ ub1 = -3.7525E-18 uc1 = -5.9821E-11 at = 1.217632E5
+ lat = -0.200775 wat = 0.128307 pat = -6.025053E-7
+ prt = 0 njs = 1.0773 xtis = 0.76
+ tpb = 1.344E-3 tpbsw = 9.9005E-4 tpbswg = 0
+ tcj = 6.7434E-4 tcjsw = 2.493E-4 tcjswg = 0
+ tvoff = 0 tvfbsdoff = 0 saref = 3E-6
+ sbref = 3E-6 wlod = 0 ku0 = -4.5E-8
+ kvsat = 0.3 kvth0 = 1.1E-8 tku0 = 0
+ llodku0 = 0 wlodku0 = 1 llodvth = 0
+ wlodvth = 1 lku0 = 0 wku0 = 2E-7
+ pku0 = 0 lkvth0 = 0 wkvth0 = 6.5E-7
+ pkvth0 = 0 stk2 = 0 lodk2 = 1
+ steta0 = 0 lodeta0 = 1

.model nhv_model.38 nmos
+ level = 54 lmin = 2E-6 lmax = 4E-6 wmin = 1E-6
+ wmax = 3E-6 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 1.16E-8
+ toxm = 1.16E-8 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 1E23 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {2.1346E-8+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {7.6507E-8-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = -4.1292E-9 dwb = -1.6944E-9 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = 0.797141 lvth0 = -9.640574E-9
+ wvth0 = 9.981546E-9 pvth0 = 4.566236E-15 k1 = 0.88325
+ k2 = -4.21037E-2 lk2 = 1.785062E-8 wk2 = 3.550394E-9
+ pk2 = -4.471189E-15 k3 = -0.884 k3b = 0.43
+ w0 = 0 lpe0 = 2.5E-8 lpeb = -2.182E-7
+ vbm = -3 dvtp0 = 0 dvtp1 = 0
+ dvt0 = 0 dvt1 = 0.53 dvt2 = -0.19251
+ dvt0w = 0.16 dvt1w = 6.9091E6 dvt2w = -0.036016
+ vfbsdoff = 0 u0 = 4.08326E-2 lu0 = 1.804126E-9
+ wu0 = -3.248109E-9 pu0 = 3.235284E-15 ua = -1.470945E-10
+ lua = -4.106334E-18 wua = -5.7213E-19 pua = 4.983634E-24
+ ub = 1.770818E-18 lub = -1.17217E-26 wub = 1.124318E-25
+ pub = -2.255559E-31 uc = 7.85112E-11 luc = -2.238024E-17
+ wuc = -3.639617E-17 puc = 6.618527E-23 ud = 0
+ up = 0 lp = 1 eu = 1.67
+ vsat = 5.366835E4 lvsat = 7.70063E-2 wvsat = 5.74254E-2
+ pvsat = -8.018068E-8 a0 = 0.66675 la0 = 8.344515E-7
+ wa0 = 4.328833E-7 pa0 = -7.992029E-13 ags = 0.191156
+ lags = -5.025416E-8 wags = -1.365754E-8 pags = 2.183093E-14
+ b0 = 3.2933E-8 b1 = 0 keta = -3.43947E-2
+ wketa = 1.202066E-8 a1 = 0 a2 = 0.659726
+ rdsw = 724.62 rdswmin = 0 rdw = 0
+ rdwmin = 0 rsw = 0 rswmin = 0
+ prwb = 0.05626 prwg = 0.048 wr = 1
+ voff = -0.20613 voffl = -4.257949E-7 minv = 0
+ nfactor = 0.946863 lnfactor = -1.85712E-7 wnfactor = 8.772754E-8
+ pnfactor = 9.564956E-14 eta0 = 0.032 etab = -0.01932
+ dsub = 0.504 cit = -8E-4 cdsc = 0
+ cdscb = 0 cdscd = 0 pclm = 0.837882
+ wpclm = 1.818103E-7 pdiblc1 = 0.21098 pdiblc2 = 2E-4
+ pdiblcb = -0.26831 drout = 0.36075 pscbe1 = 9.3731E8
+ pscbe2 = 1.68E-6 pvag = 1.99 delta = 0.0246
+ fprout = 10.125 pdits = 0 pditsl = 0
+ pditsd = 0 lambda = 0 vtl = 0
+ lc = 5E-9 xn = 3 alpha0 = 6.415903E-6
+ lalpha0 = 1.435839E-11 walpha0 = 2.051601E-11 palpha0 = -3.637902E-17
+ alpha1 = 0 beta0 = 22.318311 lbeta0 = 1.429678E-5
+ wbeta0 = 4.218632E-6 pbeta0 = -8.659755E-12 aigbacc = 1
+ bigbacc = 0 cigbacc = 0 nigbacc = 1
+ aigbinv = 0.35 bigbinv = 0.03 cigbinv = 6E-3
+ eigbinv = 1.1 nigbinv = 3 aigc = 0.43
+ bigc = 0.054 cigc = 0.075 aigsd = 0.43
+ bigsd = 0.054 cigsd = 0.075 dlcig = 0
+ nigc = 1 poxedge = 1 pigcd = 1
+ ntox = 1 toxref = 1.16E-8 agidl = 5.06E-11
+ bgidl = 1.058E9 cgidl = 4E3 egidl = 0.8
+ noia = 2.6E41 noib = 0 noic = 0
+ em = 4.1E7 af = 1 ef = 0.89
+ kf = 0 lintnoi = 0 tnoia = 7.5E6
+ tnoib = 7.2E6 ntnoi = 1 rnoia = 0.794
+ rnoib = 0.38 xpart = 0 cgso = {2.754679E-10/sw_func_tox_hv_ratio}
+ cgdo = {2.754679E-10/sw_func_tox_hv_ratio} cgbo = {0/sw_func_tox_hv_ratio} ckappas = 0.6
+ cf = 0 clc = 1E-7 cle = 0.6
+ dlc = 6.5995E-8 dwc = 0 vfbcv = -1
+ noff = 4 voffcv = -0.4104 acde = 0.4176
+ moin = 15 cgsl = {4.49025E-11/sw_func_tox_hv_ratio} cgdl = {4.49025E-11/sw_func_tox_hv_ratio}
+ ijthsrev = 0.1 ijthsfwd = 0.1 xjbvs = 1
+ bvs = 12.636 jss = 3.75E-4 jsws = 5.84E-11
+ cjs = {8.310E-04*sw_func_nsd_pw_cj} mjs = 0.295 mjsws = 0.037586
+ cjsws = {8.643094E-11*sw_func_nsd_pw_cj} cjswgs = {5.47776E-11*sw_func_nsd_pw_cj} mjswgs = 0.78692
+ pbs = 0.72468 pbsws = 0.29067 pbswgs = 0.54958
+ xrcrg1 = 12 xrcrg2 = 1 rbpb = 50
+ rbpd = 50 rbps = 50 rbdb = 50
+ rbsb = 50 gbmin = 1E-12 tnom = 30
+ ute = -1.24701 lute = -2.101265E-7 wute = 7.496672E-8
+ pute = 2.011558E-13 kt1 = -0.407353 lkt1 = 6.394796E-8
+ kt1l = 0 kt2 = -0.019151 ua1 = 3.0044E-9
+ ub1 = -3.7525E-18 uc1 = -5.9821E-11 at = 1.290087E5
+ lat = -0.228648 wat = -6.75274E-2 pat = 1.508668E-7
+ prt = 0 njs = 1.0773 xtis = 0.76
+ tpb = 1.344E-3 tpbsw = 9.9005E-4 tpbswg = 0
+ tcj = 6.7434E-4 tcjsw = 2.493E-4 tcjswg = 0
+ tvoff = 0 tvfbsdoff = 0 saref = 3E-6
+ sbref = 3E-6 wlod = 0 ku0 = -4.5E-8
+ kvsat = 0.3 kvth0 = 1.1E-8 tku0 = 0
+ llodku0 = 0 wlodku0 = 1 llodvth = 0
+ wlodvth = 1 lku0 = 0 wku0 = 2E-7
+ pku0 = 0 lkvth0 = 0 wkvth0 = 6.5E-7
+ pkvth0 = 0 stk2 = 0 lodk2 = 1
+ steta0 = 0 lodeta0 = 1

.model nhv_model.39 nmos
+ level = 54 lmin = 1E-6 lmax = 2E-6 wmin = 1E-6
+ wmax = 3E-6 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 1.16E-8
+ toxm = 1.16E-8 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 1E23 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {2.1346E-8+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {7.6507E-8-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = -4.1292E-9 dwb = -1.6944E-9 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = 0.78294 lvth0 = 1.65895E-8
+ wvth0 = 1.461189E-8 pvth0 = -3.985938E-15 k1 = 0.88325
+ k2 = -3.95294E-2 lk2 = 1.309593E-8 wk2 = 8.447246E-10
+ pk2 = 5.261439E-16 k3 = -0.884 k3b = 0.43
+ w0 = 0 lpe0 = 2.5E-8 lpeb = -2.182E-7
+ vbm = -3 dvtp0 = 0 dvtp1 = 0
+ dvt0 = 0 dvt1 = 0.53 dvt2 = -0.19251
+ dvt0w = 0.16 dvt1w = 6.9091E6 dvt2w = -0.036016
+ vfbsdoff = 0 u0 = 4.12473E-2 lu0 = 1.038092E-9
+ wu0 = -1.951289E-9 pu0 = 8.400764E-16 ua = -1.511677E-10
+ lua = 3.41687E-18 wua = 5.507302E-18 pua = -6.244991E-24
+ ub = 1.752576E-18 lub = 2.197152E-26 wub = 3.988055E-26
+ pub = -9.155479E-32 uc = 5.850306E-11 luc = 1.45745E-17
+ wuc = 2.277404E-17 puc = -4.310128E-23 ud = 0
+ up = 0 lp = 1 eu = 1.67
+ vsat = 9.313593E4 lvsat = 4.110266E-3 wvsat = 1.80901E-2
+ pvsat = -7.528995E-9 a0 = 1.118733 la0 = -3.544078E-10
+ wa0 = 2.9823E-9 pa0 = -5.18172E-15 ags = 0.159298
+ lags = 8.585532E-9 wags = 2.095676E-9 pags = -7.265037E-15
+ b0 = 3.2933E-8 b1 = 0 keta = -5.44977E-2
+ lketa = 3.712993E-8 wketa = 2.220199E-8 pketa = -1.880477E-14
+ a1 = 0 a2 = 0.659726 rdsw = 724.62
+ rdswmin = 0 rdw = 0 rdwmin = 0
+ rsw = 0 rswmin = 0 prwb = 0.05626
+ prwg = 0.048 wr = 1 voff = -0.20613
+ voffl = -4.257949E-7 minv = 0 nfactor = 0.864036
+ lnfactor = -3.273184E-8 wnfactor = 1.307142E-7 pnfactor = 1.625377E-14
+ eta0 = 0.032 etab = -0.01932 dsub = 0.504
+ cit = -8E-4 cdsc = 0 cdscb = 0
+ cdscd = 0 pclm = 0.837882 wpclm = 1.818103E-7
+ pdiblc1 = 0.21098 pdiblc2 = 2E-4 pdiblcb = -0.26831
+ drout = 0.36075 pscbe1 = 9.3731E8 pscbe2 = 1.68E-6
+ pvag = 1.99 delta = 0.0246 fprout = 10.125
+ pdits = 0 pditsl = 0 pditsd = 0
+ lambda = 0 vtl = 0 lc = 5E-9
+ xn = 3 alpha0 = 1.438483E-5 lalpha0 = -3.601001E-13
+ walpha0 = -1.062781E-11 palpha0 = 2.114319E-17 alpha1 = 0
+ beta0 = 27.317933 lbeta0 = 5.062552E-6 wbeta0 = -2.641221E-6
+ pbeta0 = 4.010297E-12 aigbacc = 1 bigbacc = 0
+ cigbacc = 0 nigbacc = 1 aigbinv = 0.35
+ bigbinv = 0.03 cigbinv = 6E-3 eigbinv = 1.1
+ nigbinv = 3 aigc = 0.43 bigc = 0.054
+ cigc = 0.075 aigsd = 0.43 bigsd = 0.054
+ cigsd = 0.075 dlcig = 0 nigc = 1
+ poxedge = 1 pigcd = 1 ntox = 1
+ toxref = 1.16E-8 agidl = 5.06E-11 bgidl = 1.058E9
+ cgidl = 4E3 egidl = 0.8 noia = 2.6E41
+ noib = 0 noic = 0 em = 4.1E7
+ af = 1 ef = 0.89 kf = 0
+ lintnoi = 0 tnoia = 7.5E6 tnoib = 7.2E6
+ ntnoi = 1 rnoia = 0.794 rnoib = 0.38
+ xpart = 0 cgso = {2.754679E-10/sw_func_tox_hv_ratio} cgdo = {2.754679E-10/sw_func_tox_hv_ratio}
+ cgbo = {0/sw_func_tox_hv_ratio} ckappas = 0.6 cf = 0
+ clc = 1E-7 cle = 0.6 dlc = 6.5995E-8
+ dwc = 0 vfbcv = -1 noff = 4
+ voffcv = -0.4104 acde = 0.4176 moin = 15
+ cgsl = {4.49025E-11/sw_func_tox_hv_ratio} cgdl = {4.49025E-11/sw_func_tox_hv_ratio} ijthsrev = 0.1
+ ijthsfwd = 0.1 xjbvs = 1 bvs = 12.636
+ jss = 3.75E-4 jsws = 5.84E-11 cjs = {8.310E-04*sw_func_nsd_pw_cj}
+ mjs = 0.295 mjsws = 0.037586 cjsws = {8.643094E-11*sw_func_nsd_pw_cj}
+ cjswgs = {5.47776E-11*sw_func_nsd_pw_cj} mjswgs = 0.78692 pbs = 0.72468
+ pbsws = 0.29067 pbswgs = 0.54958 xrcrg1 = 12
+ xrcrg2 = 1 rbpb = 50 rbpd = 50
+ rbps = 50 rbdb = 50 rbsb = 50
+ gbmin = 1E-12 tnom = 30 ute = -1.329195
+ lute = -5.833094E-8 wute = 9.048021E-8 pute = 1.725026E-13
+ kt1 = -0.37273 kt1l = 0 kt2 = -0.019151
+ ua1 = 3.0044E-9 ub1 = -3.945662E-18 lub1 = 3.567679E-25
+ wub1 = -1.801995E-25 pub1 = 3.328259E-31 uc1 = -5.9821E-11
+ at = -1.069848E4 lat = 2.93891E-2 wat = 2.61446E-2
+ pat = -2.21441E-8 prt = 0 njs = 1.0773
+ xtis = 0.76 tpb = 1.344E-3 tpbsw = 9.9005E-4
+ tpbswg = 0 tcj = 6.7434E-4 tcjsw = 2.493E-4
+ tcjswg = 0 tvoff = 0 tvfbsdoff = 0
+ saref = 3E-6 sbref = 3E-6 wlod = 0
+ ku0 = -4.5E-8 kvsat = 0.3 kvth0 = 1.1E-8
+ tku0 = 0 llodku0 = 0 wlodku0 = 1
+ llodvth = 0 wlodvth = 1 lku0 = 0
+ wku0 = 2E-7 pku0 = 0 lkvth0 = 0
+ wkvth0 = 6.5E-7 pkvth0 = 0 stk2 = 0
+ lodk2 = 1 steta0 = 0 lodeta0 = 1

.model nhv_model.40 nmos
+ level = 54 lmin = 8E-7 lmax = 1E-6 wmin = 1E-6
+ wmax = 3E-6 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 1.16E-8
+ toxm = 1.16E-8 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 1E23 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {2.1346E-8+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {7.6507E-8-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = -4.1292E-9 dwb = -1.6944E-9 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = 0.809965 lvth0 = -6.300366E-9
+ wvth0 = -1.209229E-8 pvth0 = 1.863212E-14 k1 = 0.88325
+ k2 = -1.88721E-2 lk2 = -4.400552E-9 wk2 = -1.38989E-8
+ pk2 = 1.301379E-14 k3 = -0.884 k3b = 0.43
+ w0 = 0 lpe0 = 2.5E-8 lpeb = -2.182E-7
+ vbm = -3 dvtp0 = 0 dvtp1 = 0
+ dvt0 = 0 dvt1 = 0.53 dvt2 = -0.19251
+ dvt0w = 0.16 dvt1w = 6.9091E6 dvt2w = -0.036016
+ vfbsdoff = 0 u0 = 4.26699E-2 lu0 = -1.668102E-10
+ wu0 = -1.541876E-9 pu0 = 4.933091E-16 ua = -1.394159E-10
+ lua = -6.536774E-18 wua = -2.468947E-17 pua = 1.933126E-23
+ ub = 1.931422E-18 lub = -1.29509E-25 wub = -5.204035E-25
+ pub = 3.82998E-31 uc = 1.058488E-10 luc = -2.552671E-17
+ wuc = -1.17242E-16 puc = 7.549035E-23 ud = 0
+ up = 0 lp = 1 eu = 1.67
+ vsat = 9.79327E4 lvsat = 4.74757E-5 wvsat = 9.366692E-3
+ pvsat = -1.404003E-10 a0 = 1.129403 la0 = -9.391795E-9
+ wa0 = -3.592761E-8 pa0 = 2.777443E-14 ags = 0.165697
+ lags = 3.166052E-9 wags = 4.572641E-9 pags = -9.362991E-15
+ b0 = 3.2933E-8 b1 = 0 keta = -0.01066
+ a1 = 0 a2 = 0.659726 rdsw = 724.62
+ rdswmin = 0 rdw = 0 rdwmin = 0
+ rsw = 0 rswmin = 0 prwb = 0.05626
+ prwg = 0.048 wr = 1 voff = -0.20613
+ voffl = -4.257949E-7 minv = 0 nfactor = 0.841773
+ lnfactor = -1.387549E-8 wnfactor = 1.014571E-7 pnfactor = 4.103411E-14
+ eta0 = 0.032 etab = -0.01932 dsub = 0.504
+ cit = -8E-4 cdsc = 0 cdscb = 0
+ cdscd = 0 pclm = 0.837882 wpclm = 1.818103E-7
+ pdiblc1 = 0.21098 pdiblc2 = 2E-4 pdiblcb = -0.26831
+ drout = 0.36075 pscbe1 = 9.3731E8 pscbe2 = 1.68E-6
+ pvag = 1.99 delta = 0.0246 fprout = 10.125
+ pdits = 0 pditsl = 0 pditsd = 0
+ lambda = 0 vtl = 0 lc = 5E-9
+ xn = 3 alpha0 = 1.934815E-5 lalpha0 = -4.563962E-12
+ walpha0 = -1.600333E-12 palpha0 = 1.349704E-17 alpha1 = 0
+ beta0 = 35.583624 lbeta0 = -1.938373E-6 wbeta0 = -4.674392E-6
+ pbeta0 = 5.732365E-12 aigbacc = 1 bigbacc = 0
+ cigbacc = 0 nigbacc = 1 aigbinv = 0.35
+ bigbinv = 0.03 cigbinv = 6E-3 eigbinv = 1.1
+ nigbinv = 3 aigc = 0.43 bigc = 0.054
+ cigc = 0.075 aigsd = 0.43 bigsd = 0.054
+ cigsd = 0.075 dlcig = 0 nigc = 1
+ poxedge = 1 pigcd = 1 ntox = 1
+ toxref = 1.16E-8 agidl = 5.06E-11 bgidl = 1.058E9
+ cgidl = 4E3 egidl = 0.8 noia = 2.6E41
+ noib = 0 noic = 0 em = 4.1E7
+ af = 1 ef = 0.89 kf = 0
+ lintnoi = 0 tnoia = 7.5E6 tnoib = 7.2E6
+ ntnoi = 1 rnoia = 0.794 rnoib = 0.38
+ xpart = 0 cgso = {2.754679E-10/sw_func_tox_hv_ratio} cgdo = {2.754679E-10/sw_func_tox_hv_ratio}
+ cgbo = {0/sw_func_tox_hv_ratio} ckappas = 0.6 cf = 0
+ clc = 1E-7 cle = 0.6 dlc = 6.5995E-8
+ dwc = 0 vfbcv = -1 noff = 4
+ voffcv = -0.4104 acde = 0.4176 moin = 15
+ cgsl = {4.49025E-11/sw_func_tox_hv_ratio} cgdl = {4.49025E-11/sw_func_tox_hv_ratio} ijthsrev = 0.1
+ ijthsfwd = 0.1 xjbvs = 1 bvs = 12.636
+ jss = 3.75E-4 jsws = 5.84E-11 cjs = {8.310E-04*sw_func_nsd_pw_cj}
+ mjs = 0.295 mjsws = 0.037586 cjsws = {8.643094E-11*sw_func_nsd_pw_cj}
+ cjswgs = {5.47776E-11*sw_func_nsd_pw_cj} mjswgs = 0.78692 pbs = 0.72468
+ pbsws = 0.29067 pbswgs = 0.54958 xrcrg1 = 12
+ xrcrg2 = 1 rbpb = 50 rbpd = 50
+ rbps = 50 rbdb = 50 rbsb = 50
+ gbmin = 1E-12 tnom = 30 ute = -1.640081
+ lute = 2.049849E-7 wute = 1.009865E-6 pute = -6.062034E-13
+ kt1 = -0.369633 lkt1 = -2.622967E-9 wkt1 = -9.158263E-9
+ pkt1 = 7.756921E-15 kt1l = 0 kt2 = -0.019151
+ ua1 = 1.467291E-9 lua1 = 1.30191E-15 wua1 = 4.545704E-15
+ pua1 = -3.850148E-21 ub1 = -1.200275E-18 lub1 = -1.968537E-24
+ wub1 = -6.660523E-24 pub1 = 5.821569E-30 uc1 = -5.9821E-11
+ at = 3.174206E4 lat = -6.557417E-3 wat = -2.28957E-2
+ pat = 1.93923E-8 prt = 0 njs = 1.0773
+ xtis = 0.76 tpb = 1.344E-3 tpbsw = 9.9005E-4
+ tpbswg = 0 tcj = 6.7434E-4 tcjsw = 2.493E-4
+ tcjswg = 0 tvoff = 0 tvfbsdoff = 0
+ saref = 2.81E-6 sbref = 2.81E-6 wlod = 0
+ ku0 = -4.5E-8 kvsat = 0.3 kvth0 = 1.1E-8
+ tku0 = 0 llodku0 = 0 wlodku0 = 1
+ llodvth = 0 wlodvth = 1 lku0 = 0
+ wku0 = 2E-7 pku0 = 0 lkvth0 = 0
+ wkvth0 = 6.5E-7 pkvth0 = 0 stk2 = 0
+ lodk2 = 1 steta0 = 0 lodeta0 = 1

.model nhv_model.41 nmos
+ level = 54 lmin = 6E-7 lmax = 8E-7 wmin = 1E-6
+ wmax = 3E-6 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 1.16E-8
+ toxm = 1.16E-8 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 1E23 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {2.1346E-8+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {7.6507E-8-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = -4.1292E-9 dwb = -1.6944E-9 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = 0.756365 lvth0 = 2.837814E-8
+ wvth0 = 3.1053E-8 pvth0 = -9.282273E-15 k1 = 0.88325
+ k2 = -2.27305E-2 lk2 = -1.904169E-9 wk2 = 4.814515E-9
+ pk2 = 9.064698E-16 k3 = -0.884 k3b = 0.43
+ w0 = 0 lpe0 = 2.5E-8 lpeb = -2.182E-7
+ vbm = -3 dvtp0 = 0 dvtp1 = 0
+ dvt0 = 0 dvt1 = 0.53 dvt2 = -0.19251
+ dvt0w = 0.16 dvt1w = 6.9091E6 dvt2w = -0.036016
+ vfbsdoff = 0 u0 = 3.49894E-2 lu0 = 4.802377E-9
+ wu0 = 7.547548E-10 pu0 = -9.92579E-16 ua = -1.530251E-10
+ lua = 2.268206E-18 wua = 8.599514E-18 pua = -2.206254E-24
+ ub = 5.26312E-20 lub = 1.086042E-24 wub = 8.973647E-25
+ pub = -5.342782E-31 uc = 5.945343E-11 luc = 4.490465E-18
+ wuc = 1.99635E-17 puc = -1.327969E-23 ud = 0
+ up = 0 lp = 1 eu = 1.67
+ vsat = 9.061669E4 lvsat = 4.780829E-3 wvsat = 2.46052E-2
+ pvsat = -9.999475E-9 a0 = 1.098541 la0 = 1.057519E-8
+ wa0 = 2.264884E-8 pa0 = -1.012372E-14 ags = 0.193701
+ lags = -1.495207E-8 wags = -3.202278E-8 pags = 1.431374E-14
+ b0 = 3.2933E-8 b1 = 0 keta = -0.01066
+ a1 = 0 a2 = 0.659726 rdsw = 724.62
+ rdswmin = 0 rdw = 0 rdwmin = 0
+ rsw = 0 rswmin = 0 prwb = 0.05626
+ prwg = 0.048 wr = 1 voff = -0.20613
+ voffl = -4.257949E-7 minv = 0 nfactor = 0.952023
+ lnfactor = -8.520609E-8 wnfactor = 2.729546E-8 pnfactor = 8.901567E-14
+ eta0 = 0.032 etab = -0.01932 dsub = 0.504
+ cit = -8E-4 cdsc = 0 cdscb = 0
+ cdscd = 0 pclm = 0.333814 lpclm = 3.261249E-7
+ wpclm = -8.750234E-7 ppclm = 6.837566E-13 pdiblc1 = 0.21098
+ pdiblc2 = 2E-4 pdiblcb = -0.26831 drout = 0.36075
+ pscbe1 = 9.3731E8 pscbe2 = 1.68E-6 pvag = 1.99
+ delta = 0.0246 fprout = 10.125 pdits = 0
+ pditsl = 0 pditsd = 0 lambda = 0
+ vtl = 0 lc = 5E-9 xn = 3
+ alpha0 = 5.7972E-7 lalpha0 = 7.578946E-12 walpha0 = 5.773051E-11
+ palpha0 = -2.488918E-17 alpha1 = 0 beta0 = 22.815657
+ lbeta0 = 6.322323E-6 wbeta0 = 1.354049E-5 pbeta0 = -6.052411E-12
+ aigbacc = 1 bigbacc = 0 cigbacc = 0
+ nigbacc = 1 aigbinv = 0.35 bigbinv = 0.03
+ cigbinv = 6E-3 eigbinv = 1.1 nigbinv = 3
+ aigc = 0.43 bigc = 0.054 cigc = 0.075
+ aigsd = 0.43 bigsd = 0.054 cigsd = 0.075
+ dlcig = 0 nigc = 1 poxedge = 1
+ pigcd = 1 ntox = 1 toxref = 1.16E-8
+ agidl = 5.06E-11 bgidl = 1.058E9 cgidl = 4E3
+ egidl = 0.8 noia = 2.6E41 noib = 0
+ noic = 0 em = 4.1E7 af = 1
+ ef = 0.89 kf = 0 lintnoi = 0
+ tnoia = 7.5E6 tnoib = 7.2E6 ntnoi = 1
+ rnoia = 0.794 rnoib = 0.38 xpart = 0
+ cgso = {2.754679E-10/sw_func_tox_hv_ratio} cgdo = {2.754679E-10/sw_func_tox_hv_ratio} cgbo = {0/sw_func_tox_hv_ratio}
+ ckappas = 0.6 cf = 0 clc = 1E-7
+ cle = 0.6 dlc = 6.5995E-8 dwc = 0
+ vfbcv = -1 noff = 4 voffcv = -0.4104
+ acde = 0.4176 moin = 15 cgsl = {4.49025E-11/sw_func_tox_hv_ratio}
+ cgdl = {4.49025E-11/sw_func_tox_hv_ratio} ijthsrev = 0.1 ijthsfwd = 0.1
+ xjbvs = 1 bvs = 12.636 jss = 3.75E-4
+ jsws = 5.84E-11 cjs = {8.310E-04*sw_func_nsd_pw_cj} mjs = 0.295
+ mjsws = 0.037586 cjsws = {8.643094E-11*sw_func_nsd_pw_cj} cjswgs = {5.47776E-11*sw_func_nsd_pw_cj}
+ mjswgs = 0.78692 pbs = 0.72468 pbsws = 0.29067
+ pbswgs = 0.54958 xrcrg1 = 12 xrcrg2 = 1
+ rbpb = 50 rbpd = 50 rbps = 50
+ rbdb = 50 rbsb = 50 gbmin = 1E-12
+ tnom = 30 ute = -1.377226 lute = 3.492112E-8
+ wute = 2.358253E-7 pute = -1.054106E-13 kt1 = -0.380297
+ lkt1 = 4.276174E-9 wkt1 = 9.158263E-9 pkt1 = -4.093616E-15
+ kt1l = 0 kt2 = -0.019151 ua1 = 6.760124E-9
+ lua1 = -2.122479E-15 wua1 = -4.545704E-15 pua1 = 2.031866E-21
+ ub1 = -1.065234E-17 lub1 = 4.14682E-24 wub1 = 8.473271E-24
+ pub1 = -3.969784E-30 uc1 = -5.9821E-11 at = -1.592505E4
+ lat = 2.42825E-2 wat = 2.28957E-2 pat = -1.023404E-8
+ prt = 0 njs = 1.0773 xtis = 0.76
+ tpb = 1.344E-3 tpbsw = 9.9005E-4 tpbswg = 0
+ tcj = 6.7434E-4 tcjsw = 2.493E-4 tcjswg = 0
+ tvoff = 0 tvfbsdoff = 0 saref = 2.41E-6
+ sbref = 2.41E-6 wlod = 0 ku0 = -4.5E-8
+ kvsat = 0.3 kvth0 = 1.1E-8 tku0 = 0
+ llodku0 = 0 wlodku0 = 1 llodvth = 0
+ wlodvth = 1 lku0 = 0 wku0 = 2E-7
+ pku0 = 0 lkvth0 = 0 wkvth0 = 6.5E-7
+ pkvth0 = 0 stk2 = 0 lodk2 = 1
+ steta0 = 0 lodeta0 = 1

.model nhv_model.42 nmos
+ level = 54 lmin = 5E-7 lmax = 6E-7 wmin = 1E-6
+ wmax = 3E-6 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 1.16E-8
+ toxm = 1.16E-8 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 1E23 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {2.1346E-8+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {7.6507E-8-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = -4.1292E-9 dwb = -1.6944E-9 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = 0.860205 lvth0 = -1.803681E-8
+ wvth0 = 2.002159E-8 pvth0 = -4.351388E-15 k1 = 0.88325
+ k2 = -3.924707E-3 lk2 = -1.031011E-8 wk2 = -3.334677E-9
+ pk2 = 4.549044E-15 k3 = -0.884 k3b = 0.43
+ w0 = 0 lpe0 = 2.5E-8 lpeb = -2.182E-7
+ vbm = -3 dvtp0 = 0 dvtp1 = 0
+ dvt0 = 0 dvt1 = 0.53 dvt2 = -0.19251
+ dvt0w = 0.16 dvt1w = 6.9091E6 dvt2w = -0.036016
+ vfbsdoff = 0 u0 = 3.85898E-2 lu0 = 3.193019E-9
+ wu0 = 1.036014E-9 pu0 = -1.118298E-15 ua = -1.397703E-10
+ lua = -3.656497E-18 wua = -1.950915E-17 pua = 1.035793E-23
+ ub = 7.140387E-19 lub = 7.904025E-25 wub = 4.739938E-25
+ pub = -3.450374E-31 uc = 4.794818E-11 luc = 9.633152E-18
+ wuc = 5.398807E-17 puc = -2.84882E-23 ud = 0
+ up = 0 lp = 1 eu = 1.67
+ vsat = 8.90268E4 lvsat = 5.491488E-3 wvsat = -1.98344E-2
+ pvsat = 9.864389E-9 a0 = 1.1222 ags = 0.16025
+ b0 = 3.2933E-8 b1 = 0 keta = -0.01066
+ a1 = 0 a2 = 0.659726 rdsw = 724.62
+ rdswmin = 0 rdw = 0 rdwmin = 0
+ rsw = 0 rswmin = 0 prwb = 0.05626
+ prwg = 0.048 wr = 1 voff = -0.20613
+ voffl = -4.257949E-7 minv = 0 nfactor = 0.682465
+ lnfactor = 3.528282E-8 wnfactor = 1.346917E-7 pnfactor = 4.101106E-14
+ eta0 = 0.032 etab = -0.01932 dsub = 0.504
+ cit = -8E-4 cdsc = 0 cdscb = 0
+ cdscd = 0 pclm = 0.295274 lpclm = 3.433518E-7
+ wpclm = 2.926334E-6 ppclm = -1.015397E-12 pdiblc1 = 0.21098
+ pdiblc2 = 2E-4 pdiblcb = -0.26831 drout = 0.36075
+ pscbe1 = 9.3731E8 pscbe2 = 1.68E-6 pvag = 1.99
+ delta = 0.0246 fprout = 10.125 pdits = 0
+ pditsl = 0 pditsd = 0 lambda = 0
+ vtl = 0 lc = 5E-9 xn = 3
+ alpha0 = 2.818226E-5 lalpha0 = -4.759004E-12 walpha0 = 9.155471E-12
+ palpha0 = -3.17682E-18 alpha1 = 0 beta0 = 36.96
+ aigbacc = 1 bigbacc = 0 cigbacc = 0
+ nigbacc = 1 aigbinv = 0.35 bigbinv = 0.03
+ cigbinv = 6E-3 eigbinv = 1.1 nigbinv = 3
+ aigc = 0.43 bigc = 0.054 cigc = 0.075
+ aigsd = 0.43 bigsd = 0.054 cigsd = 0.075
+ dlcig = 0 nigc = 1 poxedge = 1
+ pigcd = 1 ntox = 1 toxref = 1.16E-8
+ agidl = 5.06E-11 bgidl = 1.058E9 cgidl = 4E3
+ egidl = 0.8 noia = 2.6E41 noib = 0
+ noic = 0 em = 4.1E7 af = 1
+ ef = 0.89 kf = 0 lintnoi = 0
+ tnoia = 7.5E6 tnoib = 7.2E6 ntnoi = 1
+ rnoia = 0.794 rnoib = 0.38 xpart = 0
+ cgso = {2.754679E-10/sw_func_tox_hv_ratio} cgdo = {2.754679E-10/sw_func_tox_hv_ratio} cgbo = {0/sw_func_tox_hv_ratio}
+ ckappas = 0.6 cf = 0 clc = 1E-7
+ cle = 0.6 dlc = 6.5995E-8 dwc = 0
+ vfbcv = -1 noff = 4 voffcv = -0.4104
+ acde = 0.4176 moin = 15 cgsl = {4.49025E-11/sw_func_tox_hv_ratio}
+ cgdl = {4.49025E-11/sw_func_tox_hv_ratio} ijthsrev = 0.1 ijthsfwd = 0.1
+ xjbvs = 1 bvs = 12.636 jss = 3.75E-4
+ jsws = 5.84E-11 cjs = {8.310E-04*sw_func_nsd_pw_cj} mjs = 0.295
+ mjsws = 0.037586 cjsws = {8.643094E-11*sw_func_nsd_pw_cj} cjswgs = {5.47776E-11*sw_func_nsd_pw_cj}
+ mjswgs = 0.78692 pbs = 0.72468 pbsws = 0.29067
+ pbswgs = 0.54958 xrcrg1 = 12 xrcrg2 = 1
+ rbpb = 50 rbpd = 50 rbps = 50
+ rbdb = 50 rbsb = 50 gbmin = 1E-12
+ tnom = 30 ute = -1.042073 lute = -1.148877E-7
+ wute = -7.6524E-7 pute = 3.420516E-13 kt1 = -0.440127
+ lkt1 = 3.101958E-8 kt1l = 0 kt2 = -0.019151
+ ua1 = -1.43283E-9 lua1 = 1.539657E-15 ub1 = 9.15848E-18
+ lub1 = -4.708341E-24 wub1 = -1.063064E-23 pub1 = 4.569396E-30
+ uc1 = -5.9821E-11 at = -1.491858E4 lat = 2.38327E-2
+ wat = 4.27513E-2 pat = -1.910922E-8 prt = 0
+ njs = 1.0773 xtis = 0.76 tpb = 1.344E-3
+ tpbsw = 9.9005E-4 tpbswg = 0 tcj = 6.7434E-4
+ tcjsw = 2.493E-4 tcjswg = 0 tvoff = 0
+ tvfbsdoff = 0 saref = 2.02E-6 sbref = 2.01E-6
+ wlod = 0 ku0 = -4.5E-8 kvsat = 0.3
+ kvth0 = 1.1E-8 tku0 = 0 llodku0 = 0
+ wlodku0 = 1 llodvth = 0 wlodvth = 1
+ lku0 = 0 wku0 = 2E-7 pku0 = 0
+ lkvth0 = 0 wkvth0 = 6.5E-7 pkvth0 = 0
+ stk2 = 0 lodk2 = 1 steta0 = 0
+ lodeta0 = 1

.model nhv_model.43 nmos
+ level = 54 lmin = 8E-6 lmax = 2.02E-5 wmin = 7.5E-7
+ wmax = 1E-6 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 1.16E-8
+ toxm = 1.16E-8 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 1E23 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {2.1346E-8+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {7.6507E-8-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = -4.1292E-9 dwb = -1.6944E-9 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = 0.77701 wvth0 = 2.64561E-8
+ k1 = 0.88325 k2 = -4.93722E-2 wk2 = 1.18871E-8
+ k3 = -0.884 k3b = 0.43 w0 = 0
+ lpe0 = 2.5E-8 lpeb = -2.182E-7 vbm = -3
+ dvtp0 = 0 dvtp1 = 0 dvt0 = 0
+ dvt1 = 0.53 dvt2 = -0.19251 dvt0w = 0.16
+ dvt1w = 6.9091E6 dvt2w = -0.036016 vfbsdoff = 0
+ u0 = 3.29785E-2 wu0 = 5.337617E-9 ua = -1.573966E-10
+ wua = 8.53269E-18 ub = 1.768536E-18 wub = 1.373182E-26
+ uc = 4.032187E-11 wuc = 1.179799E-17 ud = 0
+ up = 0 lp = 1 eu = 1.67
+ vsat = 1.144463E5 wvsat = -2.437602E-3 a0 = 2.390513
+ wa0 = -1.214584E-6 ags = 0.155324 wags = 3.483875E-9
+ b0 = 5.481145E-8 wb0 = -2.094442E-14 b1 = -2.020581E-9
+ wb1 = 1.934318E-15 keta = -2.63195E-2 wketa = 4.290179E-9
+ a1 = 0 a2 = 0.659726 rdsw = 724.62
+ rdswmin = 0 rdw = 0 rdwmin = 0
+ rsw = 0 rswmin = 0 prwb = 0.05626
+ prwg = 0.048 wr = 1 voff = -0.20613
+ voffl = -4.257949E-7 minv = 0 nfactor = 1.225526
+ wnfactor = -1.356661E-7 eta0 = 0.032 etab = -0.01932
+ dsub = 0.504 cit = -8E-4 cdsc = 0
+ cdscb = 0 cdscd = 0 pclm = 3.354079
+ wpclm = -2.226966E-6 pdiblc1 = 0.21098 pdiblc2 = 2E-4
+ pdiblcb = -0.26831 drout = 0.36075 pscbe1 = 9.3731E8
+ pscbe2 = 1.68E-6 pvag = 1.99 delta = 0.0246
+ fprout = 10.125 pdits = 0 pditsl = 0
+ pditsd = 0 lambda = 0 vtl = 0
+ lc = 5E-9 xn = 3 alpha0 = 3.859256E-5
+ walpha0 = -7.445519E-12 alpha1 = 0 beta0 = 14.91913
+ wbeta0 = 1.153256E-5 aigbacc = 1 bigbacc = 0
+ cigbacc = 0 nigbacc = 1 aigbinv = 0.35
+ bigbinv = 0.03 cigbinv = 6E-3 eigbinv = 1.1
+ nigbinv = 3 aigc = 0.43 bigc = 0.054
+ cigc = 0.075 aigsd = 0.43 bigsd = 0.054
+ cigsd = 0.075 dlcig = 0 nigc = 1
+ poxedge = 1 pigcd = 1 ntox = 1
+ toxref = 1.16E-8 agidl = 5.06E-11 bgidl = 1.058E9
+ cgidl = 4E3 egidl = 0.8 noia = 2.6E41
+ noib = 0 noic = 0 em = 4.1E7
+ af = 1 ef = 0.89 kf = 0
+ lintnoi = 0 tnoia = 7.5E6 tnoib = 7.2E6
+ ntnoi = 1 rnoia = 0.794 rnoib = 0.38
+ xpart = 0 cgso = {2.754679E-10/sw_func_tox_hv_ratio} cgdo = {2.754679E-10/sw_func_tox_hv_ratio}
+ cgbo = {0/sw_func_tox_hv_ratio} ckappas = 0.6 cf = 0
+ clc = 1E-7 cle = 0.6 dlc = 6.5995E-8
+ dwc = 0 vfbcv = -1 noff = 4
+ voffcv = -0.4104 acde = 0.4176 moin = 15
+ cgsl = {4.49025E-11/sw_func_tox_hv_ratio} cgdl = {4.49025E-11/sw_func_tox_hv_ratio} ijthsrev = 0.1
+ ijthsfwd = 0.1 xjbvs = 1 bvs = 12.636
+ jss = 3.75E-4 jsws = 5.84E-11 cjs = {8.310E-04*sw_func_nsd_pw_cj}
+ mjs = 0.295 mjsws = 0.037586 cjsws = {8.643094E-11*sw_func_nsd_pw_cj}
+ cjswgs = {5.47776E-11*sw_func_nsd_pw_cj} mjswgs = 0.78692 pbs = 0.72468
+ pbsws = 0.29067 pbswgs = 0.54958 xrcrg1 = 12
+ xrcrg2 = 1 rbpb = 50 rbpd = 50
+ rbps = 50 rbdb = 50 rbsb = 50
+ gbmin = 1E-12 tnom = 30 ute = -1.1687
+ kt1 = -0.449315 wkt1 = 5.416893E-8 kt1l = 0
+ kt2 = -0.019151 ua1 = 3.0044E-9 ub1 = -3.7525E-18
+ uc1 = -5.9821E-11 at = 5.178002E5 wat = -0.352098
+ prt = 0 njs = 1.0773 xtis = 0.76
+ tpb = 1.344E-3 tpbsw = 9.9005E-4 tpbswg = 0
+ tcj = 6.7434E-4 tcjsw = 2.493E-4 tcjswg = 0
+ tvoff = 0 tvfbsdoff = 0 saref = 3E-6
+ sbref = 3E-6 wlod = 0 ku0 = -4.5E-8
+ kvsat = 0.3 kvth0 = 1.1E-8 tku0 = 0
+ llodku0 = 0 wlodku0 = 1 llodvth = 0
+ wlodvth = 1 lku0 = 0 wku0 = 2E-7
+ pku0 = 0 lkvth0 = 0 wkvth0 = 6.5E-7
+ pkvth0 = 0 stk2 = 0 lodk2 = 1
+ steta0 = 0 lodeta0 = 1

.model nhv_model.44 nmos
+ level = 54 lmin = 4E-6 lmax = 8E-6 wmin = 7.5E-7
+ wmax = 1E-6 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 1.16E-8
+ toxm = 1.16E-8 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 1E23 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {2.1346E-8+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {7.6507E-8-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = -4.1292E-9 dwb = -1.6944E-9 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = 0.770911 lvth0 = 4.78559E-8
+ wvth0 = 3.076972E-8 pvth0 = -3.384886E-14 k1 = 0.88325
+ k2 = -5.66865E-2 lk2 = 5.739529E-8 wk2 = 1.706057E-8
+ pk2 = -4.059615E-14 k3 = -0.884 k3b = 0.43
+ w0 = 0 lpe0 = 2.5E-8 lpeb = -2.182E-7
+ vbm = -3 dvtp0 = 0 dvtp1 = 0
+ dvt0 = 0 dvt1 = 0.53 dvt2 = -0.19251
+ dvt0w = 0.16 dvt1w = 6.9091E6 dvt2w = -0.036016
+ vfbsdoff = 0 u0 = 3.21207E-2 lu0 = 6.731066E-9
+ wu0 = 5.944338E-9 pu0 = -4.760936E-15 ua = -1.613633E-10
+ lua = 3.112657E-17 wua = 1.133836E-17 pua = -2.201607E-23
+ ub = 1.617212E-18 lub = 1.187439E-24 wub = 1.207647E-25
+ pub = -8.398851E-31 uc = 4.032187E-11 wuc = 1.179799E-17
+ ud = 0 up = 0 lp = 1
+ eu = 1.67 vsat = 1.144463E5 wvsat = -2.437602E-3
+ a0 = 2.401293 la0 = -8.459224E-8 wa0 = -1.222209E-6
+ pa0 = 5.983277E-14 ags = 0.115588 lags = 3.118118E-7
+ wags = 3.158983E-8 pags = -2.20547E-13 b0 = 5.481145E-8
+ wb0 = -2.094442E-14 b1 = -2.020581E-9 wb1 = 1.934318E-15
+ keta = -2.63195E-2 wketa = 4.290179E-9 a1 = 0
+ a2 = 0.659726 rdsw = 724.62 rdswmin = 0
+ rdw = 0 rdwmin = 0 rsw = 0
+ rswmin = 0 prwb = 0.05626 prwg = 0.048
+ wr = 1 voff = -0.20613 voffl = -4.257949E-7
+ minv = 0 nfactor = 1.474517 lnfactor = -1.953827E-6
+ wnfactor = -3.117792E-7 pnfactor = 1.381957E-12 eta0 = 0.032
+ etab = -0.01932 dsub = 0.504 cit = -8E-4
+ cdsc = 0 cdscb = 0 cdscd = 0
+ pclm = 3.354079 wpclm = -2.226966E-6 pdiblc1 = 0.21098
+ pdiblc2 = 2E-4 pdiblcb = -0.26831 drout = 0.36075
+ pscbe1 = 9.3731E8 pscbe2 = 1.68E-6 pvag = 1.99
+ delta = 0.0246 fprout = 10.125 pdits = 0
+ pditsl = 0 pditsd = 0 lambda = 0
+ vtl = 0 lc = 5E-9 xn = 3
+ alpha0 = 7.215715E-5 lalpha0 = -2.633809E-10 walpha0 = -3.118602E-11
+ palpha0 = 1.862914E-16 alpha1 = 0 beta0 = 10.779719
+ lbeta0 = 3.24819E-5 wbeta0 = 1.44604E-5 pbeta0 = -2.297471E-11
+ aigbacc = 1 bigbacc = 0 cigbacc = 0
+ nigbacc = 1 aigbinv = 0.35 bigbinv = 0.03
+ cigbinv = 6E-3 eigbinv = 1.1 nigbinv = 3
+ aigc = 0.43 bigc = 0.054 cigc = 0.075
+ aigsd = 0.43 bigsd = 0.054 cigsd = 0.075
+ dlcig = 0 nigc = 1 poxedge = 1
+ pigcd = 1 ntox = 1 toxref = 1.16E-8
+ agidl = 5.06E-11 bgidl = 1.058E9 cgidl = 4E3
+ egidl = 0.8 noia = 2.6E41 noib = 0
+ noic = 0 em = 4.1E7 af = 1
+ ef = 0.89 kf = 0 lintnoi = 0
+ tnoia = 7.5E6 tnoib = 7.2E6 ntnoi = 1
+ rnoia = 0.794 rnoib = 0.38 xpart = 0
+ cgso = {2.754679E-10/sw_func_tox_hv_ratio} cgdo = {2.754679E-10/sw_func_tox_hv_ratio} cgbo = {0/sw_func_tox_hv_ratio}
+ ckappas = 0.6 cf = 0 clc = 1E-7
+ cle = 0.6 dlc = 6.5995E-8 dwc = 0
+ vfbcv = -1 noff = 4 voffcv = -0.4104
+ acde = 0.4176 moin = 15 cgsl = {4.49025E-11/sw_func_tox_hv_ratio}
+ cgdl = {4.49025E-11/sw_func_tox_hv_ratio} ijthsrev = 0.1 ijthsfwd = 0.1
+ xjbvs = 1 bvs = 12.636 jss = 3.75E-4
+ jsws = 5.84E-11 cjs = {8.310E-04*sw_func_nsd_pw_cj} mjs = 0.295
+ mjsws = 0.037586 cjsws = {8.643094E-11*sw_func_nsd_pw_cj} cjswgs = {5.47776E-11*sw_func_nsd_pw_cj}
+ mjswgs = 0.78692 pbs = 0.72468 pbsws = 0.29067
+ pbswgs = 0.54958 xrcrg1 = 12 xrcrg2 = 1
+ rbpb = 50 rbpd = 50 rbps = 50
+ rbdb = 50 rbsb = 50 gbmin = 1E-12
+ tnom = 30 ute = -1.1687 kt1 = -0.45668
+ lkt1 = 5.779698E-8 wkt1 = 5.937861E-8 pkt1 = -4.088027E-14
+ kt1l = 0 kt2 = -0.019151 ua1 = 3.0044E-9
+ ub1 = -3.7525E-18 uc1 = -5.9821E-11 at = 9.229027E5
+ lat = -3.178834 wat = -0.63863 pat = 2.248415E-6
+ prt = 0 njs = 1.0773 xtis = 0.76
+ tpb = 1.344E-3 tpbsw = 9.9005E-4 tpbswg = 0
+ tcj = 6.7434E-4 tcjsw = 2.493E-4 tcjswg = 0
+ tvoff = 0 tvfbsdoff = 0 saref = 3E-6
+ sbref = 3E-6 wlod = 0 ku0 = -4.5E-8
+ kvsat = 0.3 kvth0 = 1.1E-8 tku0 = 0
+ llodku0 = 0 wlodku0 = 1 llodvth = 0
+ wlodvth = 1 lku0 = 0 wku0 = 2E-7
+ pku0 = 0 lkvth0 = 0 wkvth0 = 6.5E-7
+ pkvth0 = 0 stk2 = 0 lodk2 = 1
+ steta0 = 0 lodeta0 = 1

.model nhv_model.45 nmos
+ level = 54 lmin = 2E-6 lmax = 4E-6 wmin = 7.5E-7
+ wmax = 1E-6 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 1.16E-8
+ toxm = 1.16E-8 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 1E23 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {2.1346E-8+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {7.6507E-8-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = -4.1292E-9 dwb = -1.6944E-9 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = 0.788199 lvth0 = -1.865105E-8
+ wvth0 = 1.854173E-8 pvth0 = 1.319204E-14 k1 = 0.88325
+ k2 = -5.48862E-2 lk2 = 5.046939E-8 wk2 = 1.578717E-8
+ pk2 = -3.569741E-14 k3 = -0.884 k3b = 0.43
+ w0 = 0 lpe0 = 2.5E-8 lpeb = -2.182E-7
+ vbm = -3 dvtp0 = 0 dvtp1 = 0
+ dvt0 = 0 dvt1 = 0.53 dvt2 = -0.19251
+ dvt0w = 0.16 dvt1w = 6.9091E6 dvt2w = -0.036016
+ vfbsdoff = 0 u0 = 2.87106E-2 lu0 = 1.984955E-8
+ wu0 = 8.356307E-9 pu0 = -1.403975E-14 ua = -1.543666E-10
+ lua = 4.210431E-18 wua = 6.389553E-18 pua = -2.978071E-24
+ ub = 2.172074E-18 lub = -9.471089E-25 wub = -2.71694E-25
+ pub = 6.698977E-31 uc = -6.21897E-12 luc = 1.790419E-16
+ wuc = 4.47167E-17 puc = -1.266378E-22 ud = 0
+ up = 0 lp = 1 eu = 1.67
+ vsat = 1.211652E5 lvsat = -2.58476E-2 wvsat = -7.189941E-3
+ pvsat = 1.828218E-8 a0 = 2.379694 la0 = -1.503239E-9
+ wa0 = -1.206932E-6 pa0 = 1.063253E-15 ags = 0.223964
+ lags = -1.051111E-7 wags = -4.506576E-8 pags = 7.434594E-14
+ b0 = 5.481145E-8 wb0 = -2.094442E-14 b1 = -2.020581E-9
+ wb1 = 1.934318E-15 keta = -2.63195E-2 wketa = 4.290179E-9
+ a1 = 0 a2 = 0.659726 rdsw = 724.62
+ rdswmin = 0 rdw = 0 rdwmin = 0
+ rsw = 0 rswmin = 0 prwb = 0.05626
+ prwg = 0.048 wr = 1 voff = -0.20613
+ voffl = -4.257949E-7 minv = 0 nfactor = 1.052033
+ lnfactor = -3.28536E-7 wnfactor = -1.295275E-8 pnfactor = 2.323762E-13
+ eta0 = 0.032 etab = -0.01932 dsub = 0.504
+ cit = -8E-4 cdsc = 0 cdscb = 0
+ cdscd = 0 pclm = 3.354079 wpclm = -2.226966E-6
+ pdiblc1 = 0.21098 pdiblc2 = 2E-4 pdiblcb = -0.26831
+ drout = 0.36075 pscbe1 = 9.3731E8 pscbe2 = 1.68E-6
+ pvag = 1.99 delta = 0.0246 fprout = 10.125
+ pdits = 0 pditsl = 0 pditsd = 0
+ lambda = 0 vtl = 0 lc = 5E-9
+ xn = 3 alpha0 = 2.722681E-5 lalpha0 = -9.053447E-11
+ walpha0 = 5.935671E-13 palpha0 = 6.403575E-17 alpha1 = 0
+ beta0 = 13.996581 lbeta0 = 2.010668E-5 wbeta0 = 1.218509E-5
+ pbeta0 = -1.422161E-11 aigbacc = 1 bigbacc = 0
+ cigbacc = 0 nigbacc = 1 aigbinv = 0.35
+ bigbinv = 0.03 cigbinv = 6E-3 eigbinv = 1.1
+ nigbinv = 3 aigc = 0.43 bigc = 0.054
+ cigc = 0.075 aigsd = 0.43 bigsd = 0.054
+ cigsd = 0.075 dlcig = 0 nigc = 1
+ poxedge = 1 pigcd = 1 ntox = 1
+ toxref = 1.16E-8 agidl = 5.06E-11 bgidl = 1.058E9
+ cgidl = 4E3 egidl = 0.8 noia = 2.6E41
+ noib = 0 noic = 0 em = 4.1E7
+ af = 1 ef = 0.89 kf = 0
+ lintnoi = 0 tnoia = 7.5E6 tnoib = 7.2E6
+ ntnoi = 1 rnoia = 0.794 rnoib = 0.38
+ xpart = 0 cgso = {2.754679E-10/sw_func_tox_hv_ratio} cgdo = {2.754679E-10/sw_func_tox_hv_ratio}
+ cgbo = {0/sw_func_tox_hv_ratio} ckappas = 0.6 cf = 0
+ clc = 1E-7 cle = 0.6 dlc = 6.5995E-8
+ dwc = 0 vfbcv = -1 noff = 4
+ voffcv = -0.4104 acde = 0.4176 moin = 15
+ cgsl = {4.49025E-11/sw_func_tox_hv_ratio} cgdl = {4.49025E-11/sw_func_tox_hv_ratio} ijthsrev = 0.1
+ ijthsfwd = 0.1 xjbvs = 1 bvs = 12.636
+ jss = 3.75E-4 jsws = 5.84E-11 cjs = {8.310E-04*sw_func_nsd_pw_cj}
+ mjs = 0.295 mjsws = 0.037586 cjsws = {8.643094E-11*sw_func_nsd_pw_cj}
+ cjswgs = {5.47776E-11*sw_func_nsd_pw_cj} mjswgs = 0.78692 pbs = 0.72468
+ pbsws = 0.29067 pbswgs = 0.54958 xrcrg1 = 12
+ xrcrg2 = 1 rbpb = 50 rbpd = 50
+ rbps = 50 rbdb = 50 rbsb = 50
+ gbmin = 1E-12 tnom = 30 ute = -1.1687
+ kt1 = -0.505309 lkt1 = 2.448716E-7 wkt1 = 9.37742E-8
+ pkt1 = -1.731996E-13 kt1l = 0 kt2 = -0.019151
+ ua1 = 3.0044E-9 ub1 = -3.7525E-18 uc1 = -5.9821E-11
+ at = 1.6731E5 lat = -0.27208 wat = -0.104194
+ pat = 1.92444E-7 prt = 0 njs = 1.0773
+ xtis = 0.76 tpb = 1.344E-3 tpbsw = 9.9005E-4
+ tpbswg = 0 tcj = 6.7434E-4 tcjsw = 2.493E-4
+ tcjswg = 0 tvoff = 0 tvfbsdoff = 0
+ saref = 3E-6 sbref = 3E-6 wlod = 0
+ ku0 = -4.5E-8 kvsat = 0.3 kvth0 = 1.1E-8
+ tku0 = 0 llodku0 = 0 wlodku0 = 1
+ llodvth = 0 wlodvth = 1 lku0 = 0
+ wku0 = 2E-7 pku0 = 0 lkvth0 = 0
+ wkvth0 = 6.5E-7 pkvth0 = 0 stk2 = 0
+ lodk2 = 1 steta0 = 0 lodeta0 = 1

.model nhv_model.46 nmos
+ level = 54 lmin = 1E-6 lmax = 2E-6 wmin = 7.5E-7
+ wmax = 1E-6 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 1.16E-8
+ toxm = 1.16E-8 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 1E23 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {2.1346E-8+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {7.6507E-8-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = -4.1292E-9 dwb = -1.6944E-9 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = 0.748499 lvth0 = 5.46761E-8
+ wvth0 = 4.758288E-8 pvth0 = -4.044655E-14 k1 = 0.88325
+ k2 = -0.031081 lk2 = 6.501584E-9 wk2 = -7.242982E-9
+ pk2 = 6.838967E-15 k3 = -0.884 k3b = 0.43
+ w0 = 0 lpe0 = 2.5E-8 lpeb = -2.182E-7
+ vbm = -3 dvtp0 = 0 dvtp1 = 0
+ dvt0 = 0 dvt1 = 0.53 dvt2 = -0.19251
+ dvt0w = 0.16 dvt1w = 6.9091E6 dvt2w = -0.036016
+ vfbsdoff = 0 u0 = 3.90291E-2 lu0 = 7.914713E-10
+ wu0 = 1.722093E-10 pu0 = 1.076168E-15 ua = -1.420386E-10
+ lua = -1.855927E-17 wua = -3.232079E-18 pua = 1.479295E-23
+ ub = 1.752083E-18 lub = -1.713916E-25 wub = 4.035192E-26
+ pub = 9.355331E-32 uc = 1.538461E-10 luc = -1.16596E-16
+ wuc = -6.84986E-17 puc = 8.246928E-23 ud = 0
+ up = 0 lp = 1 eu = 1.67
+ vsat = 1.041713E5 lvsat = 5.540044E-3 wvsat = 7.52588E-3
+ pvsat = -8.897733E-9 a0 = 3.466497 la0 = -2.008813E-6
+ wa0 = -2.244552E-6 pa0 = 1.917532E-12 ags = 0.164989
+ lags = 3.815847E-9 wags = -3.351892E-9 pags = -2.698979E-15
+ b0 = -1.164185E-9 lb0 = 1.033862E-13 wb0 = 3.264151E-14
+ pb0 = -9.897245E-20 b1 = -3.366594E-9 lb1 = 2.486067E-15
+ wb1 = 3.222867E-15 pb1 = -2.379932E-21 keta = -3.95829E-2
+ lketa = 2.449728E-8 wketa = 7.923901E-9 pketa = -6.711433E-15
+ a1 = 0 a2 = 0.659726 rdsw = 724.62
+ rdswmin = 0 rdw = 0 rdwmin = 0
+ rsw = 0 rswmin = 0 prwb = 0.05626
+ prwg = 0.048 wr = 1 voff = -0.20613
+ voffl = -4.257949E-7 minv = 0 nfactor = 0.846788
+ lnfactor = 5.05478E-8 wnfactor = 1.472253E-7 pnfactor = -6.34705E-14
+ eta0 = 0.032 etab = -0.01932 dsub = 0.504
+ cit = -8E-4 cdsc = 0 cdscb = 0
+ cdscd = 0 pclm = 5.94026 lpclm = -4.776639E-6
+ wpclm = -4.702737E-6 ppclm = 4.572715E-12 pdiblc1 = 0.21098
+ pdiblc2 = 2E-4 pdiblcb = -0.26831 drout = 0.36075
+ pscbe1 = 9.3731E8 pscbe2 = 1.68E-6 pvag = 1.99
+ delta = 0.0246 fprout = 10.125 pdits = 0
+ pditsl = 0 pditsd = 0 lambda = 0
+ vtl = 0 lc = 5E-9 xn = 3
+ alpha0 = -6.683363E-5 lalpha0 = 8.319385E-11 walpha0 = 6.712327E-11
+ palpha0 = -5.884368E-17 alpha1 = 0 beta0 = 15.905411
+ lbeta0 = 1.65811E-5 wbeta0 = 8.284078E-6 pbeta0 = -7.016498E-12
+ aigbacc = 1 bigbacc = 0 cigbacc = 0
+ nigbacc = 1 aigbinv = 0.35 bigbinv = 0.03
+ cigbinv = 6E-3 eigbinv = 1.1 nigbinv = 3
+ aigc = 0.43 bigc = 0.054 cigc = 0.075
+ aigsd = 0.43 bigsd = 0.054 cigsd = 0.075
+ dlcig = 0 nigc = 1 poxedge = 1
+ pigcd = 1 ntox = 1 toxref = 1.16E-8
+ agidl = 5.06E-11 bgidl = 1.058E9 cgidl = 4E3
+ egidl = 0.8 noia = 2.6E41 noib = 0
+ noic = 0 em = 4.1E7 af = 1
+ ef = 0.89 kf = 0 lintnoi = 0
+ tnoia = 7.5E6 tnoib = 7.2E6 ntnoi = 1
+ rnoia = 0.794 rnoib = 0.38 xpart = 0
+ cgso = {2.754679E-10/sw_func_tox_hv_ratio} cgdo = {2.754679E-10/sw_func_tox_hv_ratio} cgbo = {0/sw_func_tox_hv_ratio}
+ ckappas = 0.6 cf = 0 clc = 1E-7
+ cle = 0.6 dlc = 6.5995E-8 dwc = 0
+ vfbcv = -1 noff = 4 voffcv = -0.4104
+ acde = 0.4176 moin = 15 cgsl = {4.49025E-11/sw_func_tox_hv_ratio}
+ cgdl = {4.49025E-11/sw_func_tox_hv_ratio} ijthsrev = 0.1 ijthsfwd = 0.1
+ xjbvs = 1 bvs = 12.636 jss = 3.75E-4
+ jsws = 5.84E-11 cjs = {8.310E-04*sw_func_nsd_pw_cj} mjs = 0.295
+ mjsws = 0.037586 cjsws = {8.643094E-11*sw_func_nsd_pw_cj} cjswgs = {5.47776E-11*sw_func_nsd_pw_cj}
+ mjswgs = 0.78692 pbs = 0.72468 pbsws = 0.29067
+ pbswgs = 0.54958 xrcrg1 = 12 xrcrg2 = 1
+ rbpb = 50 rbpd = 50 rbps = 50
+ rbdb = 50 rbsb = 50 gbmin = 1E-12
+ tnom = 30 ute = -1.732635 lute = 1.041581E-6
+ wute = 4.766966E-7 pute = -8.804519E-13 kt1 = -0.37273
+ kt1l = 0 kt2 = -0.019151 ua1 = 3.0044E-9
+ ub1 = -4.494065E-18 lub1 = 1.36966E-24 wub1 = 3.447906E-25
+ pub1 = -6.368235E-31 uc1 = -5.9821E-11 at = 1.661206E4
+ lat = 6.257485E-3 prt = 0 njs = 1.0773
+ xtis = 0.76 tpb = 1.344E-3 tpbsw = 9.9005E-4
+ tpbswg = 0 tcj = 6.7434E-4 tcjsw = 2.493E-4
+ tcjswg = 0 tvoff = 0 tvfbsdoff = 0
+ saref = 3E-6 sbref = 3E-6 wlod = 0
+ ku0 = -4.5E-8 kvsat = 0.3 kvth0 = 1.1E-8
+ tku0 = 0 llodku0 = 0 wlodku0 = 1
+ llodvth = 0 wlodvth = 1 lku0 = 0
+ wku0 = 2E-7 pku0 = 0 lkvth0 = 0
+ wkvth0 = 6.5E-7 pkvth0 = 0 stk2 = 0
+ lodk2 = 1 steta0 = 0 lodeta0 = 1

.model nhv_model.47 nmos
+ level = 54 lmin = 8E-7 lmax = 1E-6 wmin = 7.5E-7
+ wmax = 1E-6 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 1.16E-8
+ toxm = 1.16E-8 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 1E23 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {2.1346E-8+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {7.6507E-8-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = -4.1292E-9 dwb = -1.6944E-9 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = 0.760573 lvth0 = 4.444945E-8
+ wvth0 = 3.519133E-8 pvth0 = -2.995108E-14 k1 = 0.88325
+ k2 = -3.81123E-2 lk2 = 1.2457E-8 wk2 = 4.519966E-9
+ pk2 = -3.124085E-15 k3 = -0.884 k3b = 0.43
+ w0 = 0 lpe0 = 2.5E-8 lpeb = -2.182E-7
+ vbm = -3 dvtp0 = 0 dvtp1 = 0
+ dvt0 = 0 dvt1 = 0.53 dvt2 = -0.19251
+ dvt0w = 0.16 dvt1w = 6.9091E6 dvt2w = -0.036016
+ vfbsdoff = 0 u0 = 0.040072 lu0 = -9.187297E-11
+ wu0 = 9.450639E-10 pu0 = 4.215711E-16 ua = -2.245903E-10
+ lua = 5.136086E-17 wua = 5.684868E-17 pua = -3.609462E-23
+ ub = 1.202273E-18 lub = 2.9429E-25 wub = 1.776169E-25
+ pub = -2.27082E-32 uc = -1.970969E-10 luc = 1.806479E-16
+ wuc = 1.727704E-16 puc = -1.218822E-22 ud = 0
+ up = 0 lp = 1 eu = 1.67
+ vsat = 1.458847E5 lvsat = -2.97906E-2 wvsat = -3.65381E-2
+ pvsat = 2.842384E-8 a0 = 1.00607 la0 = 7.513436E-8
+ wa0 = 8.213954E-8 pa0 = -5.314314E-14 ags = 0.199398
+ lags = -2.532842E-8 wags = -2.768992E-8 pags = 1.791499E-14
+ b0 = 4.054649E-7 lb0 = -2.410229E-13 wb0 = -3.566278E-13
+ pb0 = 2.307332E-19 b1 = -1.826954E-9 lb1 = 1.182014E-15
+ wb1 = 1.748958E-15 pb1 = -1.131551E-21 keta = 4.59273E-2
+ lketa = -4.792861E-8 wketa = -5.417143E-8 pketa = 4.588245E-14
+ a1 = 0 a2 = 0.659726 rdsw = 724.62
+ rdswmin = 0 rdw = 0 rdwmin = 0
+ rsw = 0 rswmin = 0 prwb = 0.05626
+ prwg = 0.048 wr = 1 voff = -0.20613
+ voffl = -4.257949E-7 minv = 0 nfactor = 0.918096
+ lnfactor = -9.848585E-9 wnfactor = 2.839265E-8 pnfactor = 3.717912E-14
+ eta0 = 0.032 etab = -0.01932 dsub = 0.504
+ cit = -8E-4 cdsc = 0 cdscb = 0
+ cdscd = 0 pclm = -1.345824 lpclm = 1.394572E-6
+ wpclm = 2.272289E-6 ppclm = -1.335035E-12 pdiblc1 = 0.21098
+ pdiblc2 = 2E-4 pdiblcb = -0.26831 drout = 0.36075
+ pscbe1 = 9.3731E8 pscbe2 = 1.68E-6 pvag = 1.99
+ delta = 0.0246 fprout = 10.125 pdits = 0
+ pditsl = 0 pditsd = 0 lambda = 0
+ vtl = 0 lc = 5E-9 xn = 3
+ alpha0 = 2.699649E-5 lalpha0 = 3.721047E-12 walpha0 = -8.922157E-12
+ palpha0 = 5.565736E-18 alpha1 = 0 beta0 = 30.700773
+ lbeta0 = 4.049632E-6 aigbacc = 1 bigbacc = 0
+ cigbacc = 0 nigbacc = 1 aigbinv = 0.35
+ bigbinv = 0.03 cigbinv = 6E-3 eigbinv = 1.1
+ nigbinv = 3 aigc = 0.43 bigc = 0.054
+ cigc = 0.075 aigsd = 0.43 bigsd = 0.054
+ cigsd = 0.075 dlcig = 0 nigc = 1
+ poxedge = 1 pigcd = 1 ntox = 1
+ toxref = 1.16E-8 agidl = 5.06E-11 bgidl = 1.058E9
+ cgidl = 4E3 egidl = 0.8 noia = 2.6E41
+ noib = 0 noic = 0 em = 4.1E7
+ af = 1 ef = 0.89 kf = 0
+ lintnoi = 0 tnoia = 7.5E6 tnoib = 7.2E6
+ ntnoi = 1 rnoia = 0.794 rnoib = 0.38
+ xpart = 0 cgso = {2.754679E-10/sw_func_tox_hv_ratio} cgdo = {2.754679E-10/sw_func_tox_hv_ratio}
+ cgbo = {0/sw_func_tox_hv_ratio} ckappas = 0.6 cf = 0
+ clc = 1E-7 cle = 0.6 dlc = 6.5995E-8
+ dwc = 0 vfbcv = -1 noff = 4
+ voffcv = -0.4104 acde = 0.4176 moin = 15
+ cgsl = {4.49025E-11/sw_func_tox_hv_ratio} cgdl = {4.49025E-11/sw_func_tox_hv_ratio} ijthsrev = 0.1
+ ijthsfwd = 0.1 xjbvs = 1 bvs = 12.636
+ jss = 3.75E-4 jsws = 5.84E-11 cjs = {8.310E-04*sw_func_nsd_pw_cj}
+ mjs = 0.295 mjsws = 0.037586 cjsws = {8.643094E-11*sw_func_nsd_pw_cj}
+ cjswgs = {5.47776E-11*sw_func_nsd_pw_cj} mjswgs = 0.78692 pbs = 0.72468
+ pbsws = 0.29067 pbswgs = 0.54958 xrcrg1 = 12
+ xrcrg2 = 1 rbpb = 50 rbpd = 50
+ rbps = 50 rbdb = 50 rbsb = 50
+ gbmin = 1E-12 tnom = 30 ute = 1.904596
+ lute = -2.039103E-6 wute = -2.383483E-6 pute = 1.54208E-12
+ kt1 = -0.3792 lkt1 = 5.479881E-9 kt1l = 0
+ kt2 = -0.019151 ua1 = 6.215715E-9 lua1 = -2.719939E-15
+ ub1 = -6.356996E-18 lub1 = 2.947536E-24 wub1 = -1.723953E-24
+ pub1 = 1.115374E-30 uc1 = -5.9821E-11 at = 7.82535E3
+ lat = 1.36997E-2 prt = 0 njs = 1.0773
+ xtis = 0.76 tpb = 1.344E-3 tpbsw = 9.9005E-4
+ tpbswg = 0 tcj = 6.7434E-4 tcjsw = 2.493E-4
+ tcjswg = 0 tvoff = 0 tvfbsdoff = 0
+ saref = 2.81E-6 sbref = 2.81E-6 wlod = 0
+ ku0 = -4.5E-8 kvsat = 0.3 kvth0 = 1.1E-8
+ tku0 = 0 llodku0 = 0 wlodku0 = 1
+ llodvth = 0 wlodvth = 1 lku0 = 0
+ wku0 = 2E-7 pku0 = 0 lkvth0 = 0
+ wkvth0 = 6.5E-7 pkvth0 = 0 stk2 = 0
+ lodk2 = 1 steta0 = 0 lodeta0 = 1

.model nhv_model.48 nmos
+ level = 54 lmin = 6E-7 lmax = 8E-7 wmin = 7.5E-7
+ wmax = 1E-6 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 1.16E-8
+ toxm = 1.16E-8 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 1E23 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {2.1346E-8+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {7.6507E-8-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = -4.1292E-9 dwb = -1.6944E-9 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = 0.718705 lvth0 = 7.153738E-8
+ wvth0 = 6.710527E-8 pvth0 = -5.059896E-14 k1 = 0.88325
+ k2 = -1.31927E-2 lk2 = -3.665626E-9 wk2 = -4.316101E-9
+ pk2 = 2.592727E-15 k3 = -0.884 k3b = 0.43
+ w0 = 0 lpe0 = 2.5E-8 lpeb = -2.182E-7
+ vbm = -3 dvtp0 = 0 dvtp1 = 0
+ dvt0 = 0 dvt1 = 0.53 dvt2 = -0.19251
+ dvt0w = 0.16 dvt1w = 6.9091E6 dvt2w = -0.036016
+ vfbsdoff = 0 u0 = 1.76435E-2 lu0 = 1.44191E-8
+ wu0 = 1.736013E-8 pu0 = -1.019874E-14 ua = -1.449898E-10
+ lua = -1.395311E-19 wua = 9.072747E-19 pua = 9.869147E-26
+ ub = -1.467499E-18 lub = 2.021595E-24 wub = 2.352598E-24
+ pub = -1.429891E-30 uc = 1.376423E-10 luc = -3.592372E-17
+ wuc = -5.488728E-17 puc = 2.540914E-23 ud = 0
+ up = 0 lp = 1 eu = 1.67
+ vsat = 1.333657E5 lvsat = -0.021691 wvsat = -1.63188E-2
+ pvsat = 1.534221E-8 a0 = 1.1222 ags = 0.16025
+ b0 = 3.2933E-8 b1 = 0 keta = -2.81526E-2
+ wketa = 1.674578E-8 a1 = 0 a2 = 0.659726
+ rdsw = 724.62 rdswmin = 0 rdw = 0
+ rdwmin = 0 rsw = 0 rswmin = 0
+ prwb = 0.05626 prwg = 0.048 wr = 1
+ voff = -0.20613 voffl = -4.257949E-7 minv = 0
+ nfactor = 0.856831 lnfactor = 2.978878E-8 wnfactor = 1.184239E-7
+ pnfactor = -2.106984E-14 eta0 = 0.032 etab = -0.01932
+ dsub = 0.504 cit = -8E-4 cdsc = 0
+ cdscb = 0 cdscd = 0 pclm = -5.347862
+ lpclm = 3.983834E-6 wpclm = 4.56409E-6 ppclm = -2.817798E-12
+ pdiblc1 = 0.21098 pdiblc2 = 2E-4 pdiblcb = -0.26831
+ drout = 0.36075 pscbe1 = 9.3731E8 pscbe2 = 1.68E-6
+ pvag = 1.99 delta = 0.0246 fprout = 10.125
+ pdits = 0 pditsl = 0 pditsd = 0
+ lambda = 0 vtl = 0 lc = 5E-9
+ xn = 3 alpha0 = 1.41769E-4 lalpha0 = -7.053519E-11
+ walpha0 = -7.743116E-11 palpha0 = 4.98901E-17 alpha1 = 0
+ beta0 = 36.96 aigbacc = 1 bigbacc = 0
+ cigbacc = 0 nigbacc = 1 aigbinv = 0.35
+ bigbinv = 0.03 cigbinv = 6E-3 eigbinv = 1.1
+ nigbinv = 3 aigc = 0.43 bigc = 0.054
+ cigc = 0.075 aigsd = 0.43 bigsd = 0.054
+ cigsd = 0.075 dlcig = 0 nigc = 1
+ poxedge = 1 pigcd = 1 ntox = 1
+ toxref = 1.16E-8 agidl = 5.06E-11 bgidl = 1.058E9
+ cgidl = 4E3 egidl = 0.8 noia = 2.6E41
+ noib = 0 noic = 0 em = 4.1E7
+ af = 1 ef = 0.89 kf = 0
+ lintnoi = 0 tnoia = 7.5E6 tnoib = 7.2E6
+ ntnoi = 1 rnoia = 0.794 rnoib = 0.38
+ xpart = 0 cgso = {2.754679E-10/sw_func_tox_hv_ratio} cgdo = {2.754679E-10/sw_func_tox_hv_ratio}
+ cgbo = {0/sw_func_tox_hv_ratio} ckappas = 0.6 cf = 0
+ clc = 1E-7 cle = 0.6 dlc = 6.5995E-8
+ dwc = 0 vfbcv = -1 noff = 4
+ voffcv = -0.4104 acde = 0.4176 moin = 15
+ cgsl = {4.49025E-11/sw_func_tox_hv_ratio} cgdl = {4.49025E-11/sw_func_tox_hv_ratio} ijthsrev = 0.1
+ ijthsfwd = 0.1 xjbvs = 1 bvs = 12.636
+ jss = 3.75E-4 jsws = 5.84E-11 cjs = {8.310E-04*sw_func_nsd_pw_cj}
+ mjs = 0.295 mjsws = 0.037586 cjsws = {8.643094E-11*sw_func_nsd_pw_cj}
+ cjswgs = {5.47776E-11*sw_func_nsd_pw_cj} mjswgs = 0.78692 pbs = 0.72468
+ pbsws = 0.29067 pbswgs = 0.54958 xrcrg1 = 12
+ xrcrg2 = 1 rbpb = 50 rbpd = 50
+ rbps = 50 rbdb = 50 rbsb = 50
+ gbmin = 1E-12 tnom = 30 ute = -0.802081
+ lute = -2.879213E-7 wute = -3.147658E-7 pute = 2.036491E-13
+ kt1 = -0.37073 kt1l = 0 kt2 = -0.019151
+ ua1 = 2.0117E-9 ub1 = -1.8012E-18 uc1 = -5.9821E-11
+ at = -5.144582E4 lat = 5.20473E-2 wat = 0.0569
+ pat = -3.681348E-8 prt = 0 njs = 1.0773
+ xtis = 0.76 tpb = 1.344E-3 tpbsw = 9.9005E-4
+ tpbswg = 0 tcj = 6.7434E-4 tcjsw = 2.493E-4
+ tcjswg = 0 tvoff = 0 tvfbsdoff = 0
+ saref = 2.41E-6 sbref = 2.41E-6 wlod = 0
+ ku0 = -4.5E-8 kvsat = 0.3 kvth0 = 1.1E-8
+ tku0 = 0 llodku0 = 0 wlodku0 = 1
+ llodvth = 0 wlodvth = 1 lku0 = 0
+ wku0 = 2E-7 pku0 = 0 lkvth0 = 0
+ wkvth0 = 6.5E-7 pkvth0 = 0 stk2 = 0
+ lodk2 = 1 steta0 = 0 lodeta0 = 1

.model nhv_model.49 nmos
+ level = 54 lmin = 5E-7 lmax = 6E-7 wmin = 7.5E-7
+ wmax = 1E-6 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 1.16E-8
+ toxm = 1.16E-8 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 1E23 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {2.1346E-8+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {7.6507E-8-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = -4.1292E-9 dwb = -1.6944E-9 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = 1.050285 lvth0 = -7.66741E-8
+ wvth0 = -1.619433E-7 pvth0 = 5.178256E-14 k1 = 0.88325
+ k2 = 1.19837E-2 lk2 = -1.491915E-8 wk2 = -1.856396E-8
+ pk2 = 8.961319E-15 k3 = -0.884 k3b = 0.43
+ w0 = 0 lpe0 = 2.5E-8 lpeb = -2.182E-7
+ vbm = -3 dvtp0 = 0 dvtp1 = 0
+ dvt0 = 0 dvt1 = 0.53 dvt2 = -0.19251
+ dvt0w = 0.16 dvt1w = 6.9091E6 dvt2w = -0.036016
+ vfbsdoff = 0 u0 = 6.22063E-2 lu0 = -5.499872E-9
+ wu0 = -2.157224E-8 pu0 = 7.203476E-15 ua = -1.46617E-10
+ lua = 5.878145E-19 wua = -1.295473E-17 pua = 6.294814E-24
+ ub = 5.980236E-18 lub = -1.307438E-24 wub = -4.567379E-24
+ pub = 1.663242E-30 uc = 1.330691E-11 luc = 1.965243E-17
+ wuc = 8.715044E-17 puc = -3.807974E-23 ud = 0
+ up = 0 lp = 1 eu = 1.67
+ vsat = 7.816825E3 lvsat = 3.44276E-2 wvsat = 5.79085E-2
+ pvsat = -1.783636E-8 a0 = 1.1222 ags = 0.16025
+ b0 = 3.2933E-8 b1 = 0 keta = -8.88494E-2
+ lketa = 2.713061E-8 wketa = 7.48513E-8 pketa = -2.597235E-14
+ a1 = 0 a2 = 0.659726 rdsw = 724.62
+ rdswmin = 0 rdw = 0 rdwmin = 0
+ rsw = 0 rswmin = 0 prwb = 0.05626
+ prwg = 0.048 wr = 1 voff = -0.20613
+ voffl = -4.257949E-7 minv = 0 nfactor = 0.682629
+ lnfactor = 1.076546E-7 wnfactor = 1.345344E-7 pnfactor = -2.8271E-14
+ eta0 = 0.032 etab = -0.01932 dsub = 0.504
+ cit = -8E-4 cdsc = 0 cdscb = 0
+ cdscd = 0 pclm = 11.476075 lpclm = -3.53623E-6
+ wpclm = -7.777136E-6 ppclm = 2.698557E-12 pdiblc1 = 0.21098
+ pdiblc2 = 2E-4 pdiblcb = -0.26831 drout = 0.36075
+ pscbe1 = 9.3731E8 pscbe2 = 1.68E-6 pvag = 1.99
+ delta = 0.0246 fprout = 10.125 pdits = 0
+ pditsl = 0 pditsd = 0 lambda = 0
+ vtl = 0 lc = 5E-9 xn = 3
+ alpha0 = -1.218626E-4 lalpha0 = 4.730445E-11 walpha0 = 1.527946E-10
+ palpha0 = -5.301758E-17 alpha1 = 0 beta0 = 36.96
+ aigbacc = 1 bigbacc = 0 cigbacc = 0
+ nigbacc = 1 aigbinv = 0.35 bigbinv = 0.03
+ cigbinv = 6E-3 eigbinv = 1.1 nigbinv = 3
+ aigc = 0.43 bigc = 0.054 cigc = 0.075
+ aigsd = 0.43 bigsd = 0.054 cigsd = 0.075
+ dlcig = 0 nigc = 1 poxedge = 1
+ pigcd = 1 ntox = 1 toxref = 1.16E-8
+ agidl = 5.06E-11 bgidl = 1.058E9 cgidl = 4E3
+ egidl = 0.8 noia = 2.6E41 noib = 0
+ noic = 0 em = 4.1E7 af = 1
+ ef = 0.89 kf = 0 lintnoi = 0
+ tnoia = 7.5E6 tnoib = 7.2E6 ntnoi = 1
+ rnoia = 0.794 rnoib = 0.38 xpart = 0
+ cgso = {2.754679E-10/sw_func_tox_hv_ratio} cgdo = {2.754679E-10/sw_func_tox_hv_ratio} cgbo = {0/sw_func_tox_hv_ratio}
+ ckappas = 0.6 cf = 0 clc = 1E-7
+ cle = 0.6 dlc = 6.5995E-8 dwc = 0
+ vfbcv = -1 noff = 4 voffcv = -0.4104
+ acde = 0.4176 moin = 15 cgsl = {4.49025E-11/sw_func_tox_hv_ratio}
+ cgdl = {4.49025E-11/sw_func_tox_hv_ratio} ijthsrev = 0.1 ijthsfwd = 0.1
+ xjbvs = 1 bvs = 12.636 jss = 3.75E-4
+ jsws = 5.84E-11 cjs = {8.310E-04*sw_func_nsd_pw_cj} mjs = 0.295
+ mjsws = 0.037586 cjsws = {8.643094E-11*sw_func_nsd_pw_cj} cjswgs = {5.47776E-11*sw_func_nsd_pw_cj}
+ mjswgs = 0.78692 pbs = 0.72468 pbsws = 0.29067
+ pbswgs = 0.54958 xrcrg1 = 12 xrcrg2 = 1
+ rbpb = 50 rbpd = 50 rbps = 50
+ rbdb = 50 rbsb = 50 gbmin = 1E-12
+ tnom = 30 ute = -2.499045 lute = 4.705981E-7
+ wute = 6.295316E-7 pute = -2.184386E-13 kt1 = -0.440127
+ lkt1 = 3.101958E-8 kt1l = 0 kt2 = -0.019151
+ ua1 = -1.43283E-9 lua1 = 1.539657E-15 ub1 = -4.301348E-18
+ lub1 = 1.117531E-24 wub1 = 2.254563E-24 pub1 = -1.007758E-30
+ uc1 = -5.9821E-11 at = 1.486142E5 lat = -3.73767E-2
+ wat = -0.1138 pat = 3.948699E-8 prt = 0
+ njs = 1.0773 xtis = 0.76 tpb = 1.344E-3
+ tpbsw = 9.9005E-4 tpbswg = 0 tcj = 6.7434E-4
+ tcjsw = 2.493E-4 tcjswg = 0 tvoff = 0
+ tvfbsdoff = 0 saref = 2.41E-6 sbref = 2.41E-6
+ wlod = 0 ku0 = -4.5E-8 kvsat = 0.3
+ kvth0 = 1.1E-8 tku0 = 0 llodku0 = 0
+ wlodku0 = 1 llodvth = 0 wlodvth = 1
+ lku0 = 0 wku0 = 2E-7 pku0 = 0
+ lkvth0 = 0 wkvth0 = 6.5E-7 pkvth0 = 0
+ stk2 = 0 lodk2 = 1 steta0 = 0
+ lodeta0 = 1

.model nhv_model.50 nmos
+ level = 54 lmin = 8E-6 lmax = 2.02E-5 wmin = 4.2E-7
+ wmax = 7.5E-7 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 1.16E-8
+ toxm = 1.16E-8 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 1E23 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {2.1346E-8+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {7.6507E-8-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = -4.1292E-9 dwb = -1.6944E-9 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = 0.823428 wvth0 = -6.375838E-9
+ k1 = 0.88325 k2 = -2.46694E-2 wk2 = -5.585409E-9
+ k3 = -0.884 k3b = 0.43 w0 = 0
+ lpe0 = 2.5E-8 lpeb = -2.182E-7 vbm = -3
+ dvtp0 = 0 dvtp1 = 0 dvt0 = 0
+ dvt1 = 0.53 dvt2 = -0.19251 dvt0w = 0.16
+ dvt1w = 6.9091E6 dvt2w = -0.036016 vfbsdoff = 0
+ u0 = 3.93442E-2 wu0 = 8.35094E-10 ua = -3.212457E-10
+ wua = 1.244244E-16 ub = 1.636762E-18 wub = 1.069368E-25
+ uc = 3.285772E-11 wuc = 1.707744E-17 ud = 0
+ up = 0 lp = 1 eu = 1.67
+ vsat = 9.076257E4 wvsat = 1.43141E-2 a0 = 0.408496
+ wa0 = 1.873125E-7 ags = 0.16025 b0 = 1.446639E-8
+ wb0 = 7.59197E-15 b1 = 1.133907E-9 wb1 = -2.96876E-16
+ keta = -0.026387 wketa = 4.337899E-9 a1 = 0
+ a2 = 0.659726 rdsw = 724.62 rdswmin = 0
+ rdw = 0 rdwmin = 0 rsw = 0
+ rswmin = 0 prwb = 0.05626 prwg = 0.048
+ wr = 1 voff = -0.20613 voffl = -4.257949E-7
+ minv = 0 nfactor = 0.889291 wnfactor = 1.021557E-7
+ eta0 = 0.032 etab = -0.01932 dsub = 0.504
+ cit = -8E-4 cdsc = 0 cdscb = 0
+ cdscd = 0 pclm = -0.131034 wpclm = 2.38083E-7
+ pdiblc1 = 0.21098 pdiblc2 = 2E-4 pdiblcb = -0.26831
+ drout = 0.36075 pscbe1 = 9.3731E8 pscbe2 = 1.68E-6
+ pvag = 1.99 delta = 0.0246 fprout = 10.125
+ pdits = 0 pditsl = 0 pditsd = 0
+ lambda = 0 vtl = 0 lc = 5E-9
+ xn = 3 alpha0 = 3.638507E-5 walpha0 = -5.884145E-12
+ alpha1 = 0 beta0 = 38.021261 wbeta0 = -4.807757E-6
+ aigbacc = 1 bigbacc = 0 cigbacc = 0
+ nigbacc = 1 aigbinv = 0.35 bigbinv = 0.03
+ cigbinv = 6E-3 eigbinv = 1.1 nigbinv = 3
+ aigc = 0.43 bigc = 0.054 cigc = 0.075
+ aigsd = 0.43 bigsd = 0.054 cigsd = 0.075
+ dlcig = 0 nigc = 1 poxedge = 1
+ pigcd = 1 ntox = 1 toxref = 1.16E-8
+ agidl = 5.06E-11 bgidl = 1.058E9 cgidl = 4E3
+ egidl = 0.8 noia = 2.6E41 noib = 0
+ noic = 0 em = 4.1E7 af = 1
+ ef = 0.89 kf = 0 lintnoi = 0
+ tnoia = 7.5E6 tnoib = 7.2E6 ntnoi = 1
+ rnoia = 0.794 rnoib = 0.38 xpart = 0
+ cgso = {2.754679E-10/sw_func_tox_hv_ratio} cgdo = {2.754679E-10/sw_func_tox_hv_ratio} cgbo = {0/sw_func_tox_hv_ratio}
+ ckappas = 0.6 cf = 0 clc = 1E-7
+ cle = 0.6 dlc = 6.5995E-8 dwc = 0
+ vfbcv = -1 noff = 4 voffcv = -0.4104
+ acde = 0.4176 moin = 15 cgsl = {4.49025E-11/sw_func_tox_hv_ratio}
+ cgdl = {4.49025E-11/sw_func_tox_hv_ratio} ijthsrev = 0.1 ijthsfwd = 0.1
+ xjbvs = 1 bvs = 12.636 jss = 3.75E-4
+ jsws = 5.84E-11 cjs = {8.310E-04*sw_func_nsd_pw_cj} mjs = 0.295
+ mjsws = 0.037586 cjsws = {8.643094E-11*sw_func_nsd_pw_cj} cjswgs = {5.47776E-11*sw_func_nsd_pw_cj}
+ mjswgs = 0.78692 pbs = 0.72468 pbsws = 0.29067
+ pbswgs = 0.54958 xrcrg1 = 12 xrcrg2 = 1
+ rbpb = 50 rbpd = 50 rbps = 50
+ rbdb = 50 rbsb = 50 gbmin = 1E-12
+ tnom = 30 ute = -1.22804 wute = 4.197184E-8
+ kt1 = -0.338429 wkt1 = -2.426118E-8 kt1l = 0
+ kt2 = -0.019151 ua1 = 3.0044E-9 ub1 = -3.7525E-18
+ uc1 = -5.9821E-11 at = -1.766575E5 wat = 0.139097
+ prt = 0 njs = 1.0773 xtis = 0.76
+ tpb = 1.344E-3 tpbsw = 9.9005E-4 tpbswg = 0
+ tcj = 6.7434E-4 tcjsw = 2.493E-4 tcjswg = 0
+ tvoff = 0 tvfbsdoff = 0 saref = 3E-6
+ sbref = 3E-6 wlod = 0 ku0 = -4.5E-8
+ kvsat = 0.3 kvth0 = 1.1E-8 tku0 = 0
+ llodku0 = 0 wlodku0 = 1 llodvth = 0
+ wlodvth = 1 lku0 = 0 wku0 = 2E-7
+ pku0 = 0 lkvth0 = 0 wkvth0 = 6.5E-7
+ pkvth0 = 0 stk2 = 0 lodk2 = 1
+ steta0 = 0 lodeta0 = 1

.model nhv_model.51 nmos
+ level = 54 lmin = 4E-6 lmax = 8E-6 wmin = 4.2E-7
+ wmax = 7.5E-7 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 1.16E-8
+ toxm = 1.16E-8 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 1E23 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {2.1346E-8+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {7.6507E-8-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = -4.1292E-9 dwb = -1.6944E-9 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = 0.825162 lvth0 = -1.360747E-8
+ wvth0 = -7.602381E-9 pvth0 = 9.62467E-15 k1 = 0.88325
+ k2 = -2.16013E-2 lk2 = -2.407495E-8 wk2 = -7.755465E-9
+ pk2 = 1.70284E-14 k3 = -0.884 k3b = 0.43
+ w0 = 0 lpe0 = 2.5E-8 lpeb = -2.182E-7
+ vbm = -3 dvtp0 = 0 dvtp1 = 0
+ dvt0 = 0 dvt1 = 0.53 dvt2 = -0.19251
+ dvt0w = 0.16 dvt1w = 6.9091E6 dvt2w = -0.036016
+ vfbsdoff = 0 u0 = 0.039618 lu0 = -2.148547E-9
+ wu0 = 6.414293E-10 pu0 = 1.519685E-15 ua = -3.207628E-10
+ lua = -3.788864E-18 wua = 1.240829E-16 pua = 2.679894E-24
+ ub = 1.612424E-18 lub = 1.909791E-25 wub = 1.241512E-25
+ pub = -1.35081E-31 uc = 5.792767E-12 luc = 2.123783E-16
+ wuc = 3.62207E-17 puc = -1.502169E-22 ud = 0
+ up = 0 lp = 1 eu = 1.67
+ vsat = 8.416485E4 lvsat = 5.17722E-2 wvsat = 1.89807E-2
+ pvsat = -3.661891E-8 a0 = 0.408496 wa0 = 1.873125E-7
+ ags = 0.16025 b0 = -5.455211E-9 lb0 = 1.563245E-13
+ wb0 = 2.168268E-14 pb0 = -1.105696E-19 b1 = 7.218283E-10
+ lb1 = 3.233572E-15 wb1 = -5.409714E-18 pb1 = -2.287132E-21
+ keta = -3.27538E-2 lketa = 4.99602E-8 wketa = 8.841188E-9
+ pketa = -3.533725E-14 a1 = 0 a2 = 0.659726
+ rdsw = 724.62 rdswmin = 0 rdw = 0
+ rdwmin = 0 rsw = 0 rswmin = 0
+ prwb = 0.05626 prwg = 0.048 wr = 1
+ voff = -0.20613 voffl = -4.257949E-7 minv = 0
+ nfactor = 0.808271 lnfactor = 6.357629E-7 wnfactor = 1.594618E-7
+ pnfactor = -4.496802E-13 eta0 = 0.032 etab = -0.01932
+ dsub = 0.504 cit = -8E-4 cdsc = 0
+ cdscb = 0 cdscd = 0 pclm = -0.131034
+ wpclm = 2.38083E-7 pdiblc1 = 0.21098 pdiblc2 = 2E-4
+ pdiblcb = -0.26831 drout = 0.36075 pscbe1 = 9.3731E8
+ pscbe2 = 1.68E-6 pvag = 1.99 delta = 0.0246
+ fprout = 10.125 pdits = 0 pditsl = 0
+ pditsd = 0 lambda = 0 vtl = 0
+ lc = 5E-9 xn = 3 alpha0 = 2.962351E-5
+ lalpha0 = 5.30579E-11 walpha0 = -1.101636E-12 palpha0 = -3.752828E-17
+ alpha1 = 0 beta0 = 39.179161 lbeta0 = -9.086025E-6
+ wbeta0 = -5.626749E-6 pbeta0 = 6.426618E-12 aigbacc = 1
+ bigbacc = 0 cigbacc = 0 nigbacc = 1
+ aigbinv = 0.35 bigbinv = 0.03 cigbinv = 6E-3
+ eigbinv = 1.1 nigbinv = 3 aigc = 0.43
+ bigc = 0.054 cigc = 0.075 aigsd = 0.43
+ bigsd = 0.054 cigsd = 0.075 dlcig = 0
+ nigc = 1 poxedge = 1 pigcd = 1
+ ntox = 1 toxref = 1.16E-8 agidl = 5.06E-11
+ bgidl = 1.058E9 cgidl = 4E3 egidl = 0.8
+ noia = 2.6E41 noib = 0 noic = 0
+ em = 4.1E7 af = 1 ef = 0.89
+ kf = 0 lintnoi = 0 tnoia = 7.5E6
+ tnoib = 7.2E6 ntnoi = 1 rnoia = 0.794
+ rnoib = 0.38 xpart = 0 cgso = {2.754679E-10/sw_func_tox_hv_ratio}
+ cgdo = {2.754679E-10/sw_func_tox_hv_ratio} cgbo = {0/sw_func_tox_hv_ratio} ckappas = 0.6
+ cf = 0 clc = 1E-7 cle = 0.6
+ dlc = 6.5995E-8 dwc = 0 vfbcv = -1
+ noff = 4 voffcv = -0.4104 acde = 0.4176
+ moin = 15 cgsl = {4.49025E-11/sw_func_tox_hv_ratio} cgdl = {4.49025E-11/sw_func_tox_hv_ratio}
+ ijthsrev = 0.1 ijthsfwd = 0.1 xjbvs = 1
+ bvs = 12.636 jss = 3.75E-4 jsws = 5.84E-11
+ cjs = {8.310E-04*sw_func_nsd_pw_cj} mjs = 0.295 mjsws = 0.037586
+ cjsws = {8.643094E-11*sw_func_nsd_pw_cj} cjswgs = {5.47776E-11*sw_func_nsd_pw_cj} mjswgs = 0.78692
+ pbs = 0.72468 pbsws = 0.29067 pbswgs = 0.54958
+ xrcrg1 = 12 xrcrg2 = 1 rbpb = 50
+ rbpd = 50 rbps = 50 rbdb = 50
+ rbsb = 50 gbmin = 1E-12 tnom = 30
+ ute = -1.245524 lute = 1.371964E-7 wute = 5.433838E-8
+ pute = -9.704011E-14 kt1 = -0.325234 lkt1 = -1.035444E-7
+ wkt1 = -3.359442E-8 pkt1 = 7.323782E-14 kt1l = 0
+ kt2 = -0.019151 ua1 = 3.0044E-9 ub1 = -3.7525E-18
+ uc1 = -5.9821E-11 at = -2.99815E5 lat = 0.966415
+ wat = 0.226208 pat = -6.835529E-7 prt = 0
+ njs = 1.0773 xtis = 0.76 tpb = 1.344E-3
+ tpbsw = 9.9005E-4 tpbswg = 0 tcj = 6.7434E-4
+ tcjsw = 2.493E-4 tcjswg = 0 tvoff = 0
+ tvfbsdoff = 0 saref = 3E-6 sbref = 3E-6
+ wlod = 0 ku0 = -4.5E-8 kvsat = 0.3
+ kvth0 = 1.1E-8 tku0 = 0 llodku0 = 0
+ wlodku0 = 1 llodvth = 0 wlodvth = 1
+ lku0 = 0 wku0 = 2E-7 pku0 = 0
+ lkvth0 = 0 wkvth0 = 6.5E-7 pkvth0 = 0
+ stk2 = 0 lodk2 = 1 steta0 = 0
+ lodeta0 = 1

.model nhv_model.52 nmos
+ level = 54 lmin = 2E-6 lmax = 4E-6 wmin = 4.2E-7
+ wmax = 7.5E-7 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 1.16E-8
+ toxm = 1.16E-8 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 1E23 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {2.1346E-8+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {7.6507E-8-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = -4.1292E-9 dwb = -1.6944E-9 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = 0.813468 lvth0 = 3.137869E-8
+ wvth0 = 6.687864E-10 pvth0 = -2.21944E-14 k1 = 0.88325
+ k2 = -2.27076E-2 lk2 = -1.981914E-8 wk2 = -6.972992E-9
+ pk2 = 1.401824E-14 k3 = -0.884 k3b = 0.43
+ w0 = 0 lpe0 = 2.5E-8 lpeb = -2.182E-7
+ vbm = -3 dvtp0 = 0 dvtp1 = 0
+ dvt0 = 0 dvt1 = 0.53 dvt2 = -0.19251
+ dvt0w = 0.16 dvt1w = 6.9091E6 dvt2w = -0.036016
+ vfbsdoff = 0 u0 = 4.10358E-2 lu0 = -7.602782E-9
+ wu0 = -3.613879E-10 pu0 = 5.377508E-15 ua = -4.009079E-10
+ lua = 3.04528E-16 wua = 1.807701E-16 pua = -2.153951E-22
+ ub = 1.630171E-18 lub = 1.227039E-25 wub = 1.115981E-25
+ pub = -8.678943E-32 uc = 6.87029E-11 luc = -2.96361E-17
+ wuc = -8.276139E-18 puc = 2.096185E-23 ud = 0
+ up = 0 lp = 1 eu = 1.67
+ vsat = 9.551095E4 lvsat = 8.123932E-3 wvsat = 1.09555E-2
+ pvsat = -5.746122E-9 a0 = 0.306117 la0 = 3.938482E-7
+ wa0 = 2.597255E-7 pa0 = -2.78572E-13 ags = 0.16025
+ b0 = 4.063506E-8 lb0 = -2.098412E-14 wb0 = -1.091734E-14
+ pb0 = 1.484223E-20 b1 = 4.06362E-9 lb1 = -9.622253E-15
+ wb1 = -2.369086E-15 pb1 = 6.805897E-21 keta = -1.97669E-2
+ wketa = -3.445087E-10 a1 = 0 a2 = 0.659726
+ rdsw = 724.62 rdswmin = 0 rdw = 0
+ rdwmin = 0 rsw = 0 rswmin = 0
+ prwb = 0.05626 prwg = 0.048 wr = 1
+ voff = -0.20613 voffl = -4.257949E-7 minv = 0
+ nfactor = 0.910043 lnfactor = 2.44246E-7 wnfactor = 8.747743E-8
+ pnfactor = -1.727572E-13 eta0 = 0.032 etab = -0.01932
+ dsub = 0.504 cit = -8E-4 cdsc = 0
+ cdscb = 0 cdscd = 0 pclm = -0.131034
+ wpclm = 2.38083E-7 pdiblc1 = 0.21098 pdiblc2 = 2E-4
+ pdiblcb = -0.26831 drout = 0.36075 pscbe1 = 9.3731E8
+ pscbe2 = 1.68E-6 pvag = 1.99 delta = 0.0246
+ fprout = 10.125 pdits = 0 pditsl = 0
+ pditsd = 0 lambda = 0 vtl = 0
+ lc = 5E-9 xn = 3 alpha0 = 4.475971E-5
+ lalpha0 = -5.170883E-12 walpha0 = -1.18076E-11 palpha0 = 3.657407E-18
+ alpha1 = 0 beta0 = 40.60898 lbeta0 = -1.458652E-5
+ wbeta0 = -6.638072E-6 pbeta0 = 1.031716E-11 aigbacc = 1
+ bigbacc = 0 cigbacc = 0 nigbacc = 1
+ aigbinv = 0.35 bigbinv = 0.03 cigbinv = 6E-3
+ eigbinv = 1.1 nigbinv = 3 aigc = 0.43
+ bigc = 0.054 cigc = 0.075 aigsd = 0.43
+ bigsd = 0.054 cigsd = 0.075 dlcig = 0
+ nigc = 1 poxedge = 1 pigcd = 1
+ ntox = 1 toxref = 1.16E-8 agidl = 5.06E-11
+ bgidl = 1.058E9 cgidl = 4E3 egidl = 0.8
+ noia = 2.6E41 noib = 0 noic = 0
+ em = 4.1E7 af = 1 ef = 0.89
+ kf = 0 lintnoi = 0 tnoia = 7.5E6
+ tnoib = 7.2E6 ntnoi = 1 rnoia = 0.794
+ rnoib = 0.38 xpart = 0 cgso = {2.754679E-10/sw_func_tox_hv_ratio}
+ cgdo = {2.754679E-10/sw_func_tox_hv_ratio} cgbo = {0/sw_func_tox_hv_ratio} ckappas = 0.6
+ cf = 0 clc = 1E-7 cle = 0.6
+ dlc = 6.5995E-8 dwc = 0 vfbcv = -1
+ noff = 4 voffcv = -0.4104 acde = 0.4176
+ moin = 15 cgsl = {4.49025E-11/sw_func_tox_hv_ratio} cgdl = {4.49025E-11/sw_func_tox_hv_ratio}
+ ijthsrev = 0.1 ijthsfwd = 0.1 xjbvs = 1
+ bvs = 12.636 jss = 3.75E-4 jsws = 5.84E-11
+ cjs = {8.310E-04*sw_func_nsd_pw_cj} mjs = 0.295 mjsws = 0.037586
+ cjsws = {8.643094E-11*sw_func_nsd_pw_cj} cjswgs = {5.47776E-11*sw_func_nsd_pw_cj} mjswgs = 0.78692
+ pbs = 0.72468 pbsws = 0.29067 pbswgs = 0.54958
+ xrcrg1 = 12 xrcrg2 = 1 rbpb = 50
+ rbpd = 50 rbps = 50 rbdb = 50
+ rbsb = 50 gbmin = 1E-12 tnom = 30
+ ute = -1.247873 lute = 1.462308E-7 wute = 5.599945E-8
+ pute = -1.034302E-13 kt1 = -0.333144 lkt1 = -7.311539E-8
+ wkt1 = -2.799972E-8 pkt1 = 5.17151E-14 kt1l = 0
+ kt2 = -0.019151 ua1 = 3.0044E-9 ub1 = -3.7525E-18
+ uc1 = -5.9821E-11 at = -1.119544E5 lat = 0.243718
+ wat = 9.33324E-2 pat = -1.723837E-7 prt = 0
+ njs = 1.0773 xtis = 0.76 tpb = 1.344E-3
+ tpbsw = 9.9005E-4 tpbswg = 0 tcj = 6.7434E-4
+ tcjsw = 2.493E-4 tcjswg = 0 tvoff = 0
+ tvfbsdoff = 0 saref = 3E-6 sbref = 3E-6
+ wlod = 0 ku0 = -4.5E-8 kvsat = 0.3
+ kvth0 = 1.1E-8 tku0 = 0 llodku0 = 0
+ wlodku0 = 1 llodvth = 0 wlodvth = 1
+ lku0 = 0 wku0 = 2E-7 pku0 = 0
+ lkvth0 = 0 wkvth0 = 6.5E-7 pkvth0 = 0
+ stk2 = 0 lodk2 = 1 steta0 = 0
+ lodeta0 = 1

.model nhv_model.53 nmos
+ level = 54 lmin = 1E-6 lmax = 2E-6 wmin = 4.2E-7
+ wmax = 7.5E-7 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 1.16E-8
+ toxm = 1.16E-8 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 1E23 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {2.1346E-8+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {7.6507E-8-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = -4.1292E-9 dwb = -1.6944E-9 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = 0.827068 lvth0 = 6.260205E-9
+ wvth0 = -7.990075E-9 pvth0 = -6.201601E-15 k1 = 0.88325
+ k2 = -4.16777E-2 lk2 = 1.521832E-8 wk2 = 2.521259E-10
+ pk2 = 6.73548E-16 k3 = -0.884 k3b = 0.43
+ w0 = 0 lpe0 = 2.5E-8 lpeb = -2.182E-7
+ vbm = -3 dvtp0 = 0 dvtp1 = 0
+ dvt0 = 0 dvt1 = 0.53 dvt2 = -0.19251
+ dvt0w = 0.16 dvt1w = 6.9091E6 dvt2w = -0.036016
+ vfbsdoff = 0 u0 = 3.59493E-2 lu0 = 1.791994E-9
+ wu0 = 2.350608E-9 pu0 = 3.684904E-16 ua = -2.361205E-10
+ lua = 1.680172E-19 wua = 6.331279E-17 pua = 1.546984E-24
+ ub = 1.656236E-18 lub = 7.456255E-26 wub = 1.081452E-25
+ pub = -8.041206E-32 uc = 5.265724E-11 wuc = 3.073083E-18
+ ud = 0 up = 0 lp = 1
+ eu = 1.67 vsat = 1.110323E5 lvsat = -2.05439E-2
+ wvsat = 2.67298E-3 pvsat = 9.551629E-9 a0 = 8.754591E-3
+ la0 = 9.430727E-7 wa0 = 2.011374E-7 pa0 = -1.703606E-13
+ ags = 0.16025 b0 = 1.208863E-7 lb0 = -1.692071E-13
+ wb0 = -5.368578E-14 pb0 = 9.383495E-20 b1 = -1.839667E-9
+ lb1 = 1.281035E-15 wb1 = 2.142859E-15 pb1 = -1.527603E-21
+ keta = -2.74804E-2 lketa = 1.424662E-8 wketa = -6.363028E-10
+ pketa = 5.389396E-16 a1 = 0 a2 = 0.659726
+ rdsw = 724.62 rdswmin = 0 rdw = 0
+ rdwmin = 0 rsw = 0 rswmin = 0
+ prwb = 0.05626 prwg = 0.048 wr = 1
+ voff = -0.20613 voffl = -4.257949E-7 minv = 0
+ nfactor = 1.053487 lnfactor = -2.069301E-8 wnfactor = 1.025306E-9
+ pnfactor = -1.30813E-14 eta0 = 0.032 etab = -0.01932
+ dsub = 0.504 cit = -8E-4 cdsc = 0
+ cdscb = 0 cdscd = 0 pclm = -1.474035
+ lpclm = 2.480503E-6 wpclm = 5.41453E-7 ppclm = -5.6032E-13
+ pdiblc1 = 0.21098 pdiblc2 = 2E-4 pdiblcb = -0.26831
+ drout = 0.36075 pscbe1 = 9.3731E8 pscbe2 = 1.68E-6
+ pvag = 1.99 delta = 0.0246 fprout = 10.125
+ pdits = 0 pditsl = 0 pditsd = 0
+ lambda = 0 vtl = 0 lc = 5E-9
+ xn = 3 alpha0 = 4.05588E-5 lalpha0 = 2.588156E-12
+ walpha0 = -8.836254E-12 palpha0 = -1.830623E-18 alpha1 = 0
+ beta0 = 27.501358 lbeta0 = 9.623074E-6 wbeta0 = 8.217166E-8
+ pbeta0 = -2.095033E-12 aigbacc = 1 bigbacc = 0
+ cigbacc = 0 nigbacc = 1 aigbinv = 0.35
+ bigbinv = 0.03 cigbinv = 6E-3 eigbinv = 1.1
+ nigbinv = 3 aigc = 0.43 bigc = 0.054
+ cigc = 0.075 aigsd = 0.43 bigsd = 0.054
+ cigsd = 0.075 dlcig = 0 nigc = 1
+ poxedge = 1 pigcd = 1 ntox = 1
+ toxref = 1.16E-8 agidl = 5.06E-11 bgidl = 1.058E9
+ cgidl = 4E3 egidl = 0.8 noia = 2.6E41
+ noib = 0 noic = 0 em = 4.1E7
+ af = 1 ef = 0.89 kf = 0
+ lintnoi = 0 tnoia = 7.5E6 tnoib = 7.2E6
+ ntnoi = 1 rnoia = 0.794 rnoib = 0.38
+ xpart = 0 cgso = {2.754679E-10/sw_func_tox_hv_ratio} cgdo = {2.754679E-10/sw_func_tox_hv_ratio}
+ cgbo = {0/sw_func_tox_hv_ratio} ckappas = 0.6 cf = 0
+ clc = 1E-7 cle = 0.6 dlc = 6.5995E-8
+ dwc = 0 vfbcv = -1 noff = 4
+ voffcv = -0.4104 acde = 0.4176 moin = 15
+ cgsl = {4.49025E-11/sw_func_tox_hv_ratio} cgdl = {4.49025E-11/sw_func_tox_hv_ratio} ijthsrev = 0.1
+ ijthsfwd = 0.1 xjbvs = 1 bvs = 12.636
+ jss = 3.75E-4 jsws = 5.84E-11 cjs = {8.310E-04*sw_func_nsd_pw_cj}
+ mjs = 0.295 mjsws = 0.037586 cjsws = {8.643094E-11*sw_func_nsd_pw_cj}
+ cjswgs = {5.47776E-11*sw_func_nsd_pw_cj} mjswgs = 0.78692 pbs = 0.72468
+ pbsws = 0.29067 pbswgs = 0.54958 xrcrg1 = 12
+ xrcrg2 = 1 rbpb = 50 rbpd = 50
+ rbps = 50 rbdb = 50 rbsb = 50
+ gbmin = 1E-12 tnom = 30 ute = -1.058677
+ lute = -2.032118E-7 kt1 = -0.37273 kt1l = 0
+ kt2 = -0.019151 ua1 = 3.0044E-9 ub1 = -4.297118E-18
+ lub1 = 1.005902E-24 wub1 = 2.054888E-25 pub1 = -3.795349E-31
+ uc1 = -5.9821E-11 at = 1.661206E4 lat = 6.257485E-3
+ prt = 0 njs = 1.0773 xtis = 0.76
+ tpb = 1.344E-3 tpbsw = 9.9005E-4 tpbswg = 0
+ tcj = 6.7434E-4 tcjsw = 2.493E-4 tcjswg = 0
+ tvoff = 0 tvfbsdoff = 0 saref = 3E-6
+ sbref = 3E-6 wlod = 0 ku0 = -4.5E-8
+ kvsat = 0.3 kvth0 = 1.1E-8 tku0 = 0
+ llodku0 = 0 wlodku0 = 1 llodvth = 0
+ wlodvth = 1 lku0 = 0 wku0 = 2E-7
+ pku0 = 0 lkvth0 = 0 wkvth0 = 6.5E-7
+ pkvth0 = 0 stk2 = 0 lodk2 = 1
+ steta0 = 0 lodeta0 = 1

.model nhv_model.54 nmos
+ level = 54 lmin = 8E-7 lmax = 1E-6 wmin = 4.2E-7
+ wmax = 7.5E-7 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 1.16E-8
+ toxm = 1.16E-8 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 1E23 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {2.1346E-8+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {7.6507E-8-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = -4.1292E-9 dwb = -1.6944E-9 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = 0.841336 lvth0 = -5.82467E-9
+ wvth0 = -2.193341E-8 pvth0 = 5.608205E-15 k1 = 0.88325
+ k2 = -3.27907E-2 lk2 = 7.691212E-9 wk2 = 7.559731E-10
+ pk2 = 2.467965E-16 k3 = -0.884 k3b = 0.43
+ w0 = 0 lpe0 = 2.5E-8 lpeb = -2.182E-7
+ vbm = -3 dvtp0 = 0 dvtp1 = 0
+ dvt0 = 0 dvt1 = 0.53 dvt2 = -0.19251
+ dvt0w = 0.16 dvt1w = 6.9091E6 dvt2w = -0.036016
+ vfbsdoff = 0 u0 = 3.71635E-2 lu0 = 7.635392E-10
+ wu0 = 3.002282E-9 pu0 = -1.834687E-16 ua = -3.583973E-10
+ lua = 1.037348E-16 wua = 1.514914E-16 pua = -7.313911E-23
+ ub = 1.221785E-18 lub = 4.425363E-25 wub = 1.638155E-25
+ pub = -1.27564E-31 uc = 9.588275E-14 luc = 4.451873E-17
+ wuc = 3.329435E-17 puc = -2.559699E-23 ud = 0
+ up = 0 lp = 1 eu = 1.67
+ vsat = 3.921944E4 lvsat = 4.02807E-2 wvsat = 3.89071E-2
+ pvsat = -2.113813E-8 a0 = 1.1222 ags = 0.16025
+ b0 = -4.406262E-7 lb0 = 3.063861E-13 wb0 = 2.418192E-13
+ pb0 = -1.564536E-19 b1 = -1.385687E-9 lb1 = 8.965201E-16
+ wb1 = 1.436846E-15 pb1 = -9.296193E-22 keta = -5.35291E-2
+ lketa = 3.630956E-8 wketa = 1.617487E-8 pketa = -1.369989E-14
+ a1 = 0 a2 = 0.659726 rdsw = 724.62
+ rdswmin = 0 rdw = 0 rdwmin = 0
+ rsw = 0 rswmin = 0 prwb = 0.05626
+ prwg = 0.048 wr = 1 voff = -0.20613
+ voffl = -4.257949E-7 minv = 0 nfactor = 0.988647
+ lnfactor = 3.422597E-8 wnfactor = -2.150888E-8 pnfactor = 6.004835E-15
+ eta0 = 0.032 etab = -0.01932 dsub = 0.504
+ cit = -8E-4 cdsc = 0 cdscb = 0
+ cdscd = 0 pclm = 2.701945 lpclm = -1.056494E-6
+ wpclm = -5.907305E-7 ppclm = 3.986235E-13 pdiblc1 = 0.21098
+ pdiblc2 = 2E-4 pdiblcb = -0.26831 drout = 0.36075
+ pscbe1 = 9.3731E8 pscbe2 = 1.68E-6 pvag = 1.99
+ delta = 0.0246 fprout = 10.125 pdits = 0
+ pditsl = 0 pditsd = 0 lambda = 0
+ vtl = 0 lc = 5E-9 xn = 3
+ alpha0 = -2.837335E-6 lalpha0 = 3.934407E-11 walpha0 = 1.217955E-11
+ palpha0 = -1.963071E-17 alpha1 = 0 beta0 = 28.61503
+ lbeta0 = 8.679809E-6 wbeta0 = 1.475263E-6 pbeta0 = -3.274961E-12
+ aigbacc = 1 bigbacc = 0 cigbacc = 0
+ nigbacc = 1 aigbinv = 0.35 bigbinv = 0.03
+ cigbinv = 6E-3 eigbinv = 1.1 nigbinv = 3
+ aigc = 0.43 bigc = 0.054 cigc = 0.075
+ aigsd = 0.43 bigsd = 0.054 cigsd = 0.075
+ dlcig = 0 nigc = 1 poxedge = 1
+ pigcd = 1 ntox = 1 toxref = 1.16E-8
+ agidl = 5.06E-11 bgidl = 1.058E9 cgidl = 4E3
+ egidl = 0.8 noia = 2.6E41 noib = 0
+ noic = 0 em = 4.1E7 af = 1
+ ef = 0.89 kf = 0 lintnoi = 0
+ tnoia = 7.5E6 tnoib = 7.2E6 ntnoi = 1
+ rnoia = 0.794 rnoib = 0.38 xpart = 0
+ cgso = {2.754679E-10/sw_func_tox_hv_ratio} cgdo = {2.754679E-10/sw_func_tox_hv_ratio} cgbo = {0/sw_func_tox_hv_ratio}
+ ckappas = 0.6 cf = 0 clc = 1E-7
+ cle = 0.6 dlc = 6.5995E-8 dwc = 0
+ vfbcv = -1 noff = 4 voffcv = -0.4104
+ acde = 0.4176 moin = 15 cgsl = {4.49025E-11/sw_func_tox_hv_ratio}
+ cgdl = {4.49025E-11/sw_func_tox_hv_ratio} ijthsrev = 0.1 ijthsfwd = 0.1
+ xjbvs = 1 bvs = 12.636 jss = 3.75E-4
+ jsws = 5.84E-11 cjs = {8.310E-04*sw_func_nsd_pw_cj} mjs = 0.295
+ mjsws = 0.037586 cjsws = {8.643094E-11*sw_func_nsd_pw_cj} cjswgs = {5.47776E-11*sw_func_nsd_pw_cj}
+ mjswgs = 0.78692 pbs = 0.72468 pbsws = 0.29067
+ pbswgs = 0.54958 xrcrg1 = 12 xrcrg2 = 1
+ rbpb = 50 rbpd = 50 rbps = 50
+ rbdb = 50 rbsb = 50 gbmin = 1E-12
+ tnom = 30 ute = -1.465199 lute = 1.411069E-7
+ kt1 = -0.3792 lkt1 = 5.479881E-9 kt1l = 0
+ kt2 = -0.019151 ua1 = 6.215715E-9 lua1 = -2.719939E-15
+ ub1 = -7.341728E-18 lub1 = 3.584644E-24 wub1 = -1.027444E-24
+ pub1 = 6.647418E-31 uc1 = -5.9821E-11 at = 7.82535E3
+ lat = 1.36997E-2 prt = 0 njs = 1.0773
+ xtis = 0.76 tpb = 1.344E-3 tpbsw = 9.9005E-4
+ tpbswg = 0 tcj = 6.7434E-4 tcjsw = 2.493E-4
+ tcjswg = 0 tvoff = 0 tvfbsdoff = 0
+ saref = 2.81E-6 sbref = 2.81E-6 wlod = 0
+ ku0 = -4.5E-8 kvsat = 0.3 kvth0 = 1.1E-8
+ tku0 = 0 llodku0 = 0 wlodku0 = 1
+ llodvth = 0 wlodvth = 1 lku0 = 0
+ wku0 = 2E-7 pku0 = 0 lkvth0 = 0
+ wkvth0 = 6.5E-7 pkvth0 = 0 stk2 = 0
+ lodk2 = 1 steta0 = 0 lodeta0 = 1

.model nhv_model.55 nmos
+ level = 54 lmin = 6E-7 lmax = 8E-7 wmin = 4.2E-7
+ wmax = 7.5E-7 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 1.16E-8
+ toxm = 1.16E-8 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 1E23 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {2.1346E-8+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {7.6507E-8-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = -4.1292E-9 dwb = -1.6944E-9 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = 0.839726 lvth0 = -4.782878E-9
+ wvth0 = -1.849402E-8 pvth0 = 3.382968E-15 k1 = 0.88325
+ k2 = -1.04959E-2 lk2 = -6.733228E-9 wk2 = -6.223574E-9
+ pk2 = 4.762466E-15 k3 = -0.884 k3b = 0.43
+ w0 = 0 lpe0 = 2.5E-8 lpeb = -2.182E-7
+ vbm = -3 dvtp0 = 0 dvtp1 = 0
+ dvt0 = 0 dvt1 = 0.53 dvt2 = -0.19251
+ dvt0w = 0.16 dvt1w = 6.9091E6 dvt2w = -0.036016
+ vfbsdoff = 0 u0 = 4.23392E-2 lu0 = -2.585036E-9
+ wu0 = -1.073448E-10 pu0 = 1.828416E-15 ua = -1.93968E-10
+ lua = -2.648686E-18 wua = 3.554992E-17 pua = 1.873437E-24
+ ub = 2.447792E-18 lub = -3.506728E-25 wub = -4.167189E-25
+ pub = 2.480336E-31 uc = 6.890531E-11 wuc = -6.269089E-18
+ ud = 0 up = 0 lp = 1
+ eu = 1.67 vsat = 9.431503E4 lvsat = 4.634581E-3
+ wvsat = 1.13021E-2 pvsat = -3.278076E-9 a0 = 1.1222
+ ags = 0.16025 b0 = 3.2933E-8 b1 = 0
+ keta = 2.591951E-3 wketa = -5.000067E-9 a1 = 0
+ a2 = 0.659726 rdsw = 724.62 rdswmin = 0
+ rdw = 0 rdwmin = 0 rsw = 0
+ rswmin = 0 prwb = 0.05626 prwg = 0.048
+ wr = 1 voff = -0.20613 voffl = -4.257949E-7
+ minv = 0 nfactor = 0.990186 lnfactor = 3.32305E-8
+ wnfactor = 2.410113E-8 pnfactor = -2.35042E-14 eta0 = 0.032
+ etab = -0.01932 dsub = 0.504 cit = -8E-4
+ cdsc = 0 cdscb = 0 cdscd = 0
+ pclm = 2.172388 lpclm = -7.138772E-7 wpclm = -7.550425E-7
+ ppclm = 5.049311E-13 pdiblc1 = 0.21098 pdiblc2 = 2E-4
+ pdiblcb = -0.26831 drout = 0.36075 pscbe1 = 9.3731E8
+ pscbe2 = 1.68E-6 pvag = 1.99 delta = 0.0246
+ fprout = 10.125 pdits = 0 pditsl = 0
+ pditsd = 0 lambda = 0 vtl = 0
+ lc = 5E-9 xn = 3 alpha0 = 5.797398E-5
+ walpha0 = -1.816224E-11 alpha1 = 0 beta0 = 45.355268
+ lbeta0 = -2.15089E-6 wbeta0 = -5.93804E-6 pbeta0 = 1.521342E-12
+ aigbacc = 1 bigbacc = 0 cigbacc = 0
+ nigbacc = 1 aigbinv = 0.35 bigbinv = 0.03
+ cigbinv = 6E-3 eigbinv = 1.1 nigbinv = 3
+ aigc = 0.43 bigc = 0.054 cigc = 0.075
+ aigsd = 0.43 bigsd = 0.054 cigsd = 0.075
+ dlcig = 0 nigc = 1 poxedge = 1
+ pigcd = 1 ntox = 1 toxref = 1.16E-8
+ agidl = 5.06E-11 bgidl = 1.058E9 cgidl = 4E3
+ egidl = 0.8 noia = 2.6E41 noib = 0
+ noic = 0 em = 4.1E7 af = 1
+ ef = 0.89 kf = 0 lintnoi = 0
+ tnoia = 7.5E6 tnoib = 7.2E6 ntnoi = 1
+ rnoia = 0.794 rnoib = 0.38 xpart = 0
+ cgso = {2.754679E-10/sw_func_tox_hv_ratio} cgdo = {2.754679E-10/sw_func_tox_hv_ratio} cgbo = {0/sw_func_tox_hv_ratio}
+ ckappas = 0.6 cf = 0 clc = 1E-7
+ cle = 0.6 dlc = 6.5995E-8 dwc = 0
+ vfbcv = -1 noff = 4 voffcv = -0.4104
+ acde = 0.4176 moin = 15 cgsl = {4.49025E-11/sw_func_tox_hv_ratio}
+ cgdl = {4.49025E-11/sw_func_tox_hv_ratio} ijthsrev = 0.1 ijthsfwd = 0.1
+ xjbvs = 1 bvs = 12.636 jss = 3.75E-4
+ jsws = 5.84E-11 cjs = {8.310E-04*sw_func_nsd_pw_cj} mjs = 0.295
+ mjsws = 0.037586 cjsws = {8.643094E-11*sw_func_nsd_pw_cj} cjswgs = {5.47776E-11*sw_func_nsd_pw_cj}
+ mjswgs = 0.78692 pbs = 0.72468 pbsws = 0.29067
+ pbswgs = 0.54958 xrcrg1 = 12 xrcrg2 = 1
+ rbpb = 50 rbpd = 50 rbps = 50
+ rbdb = 50 rbsb = 50 gbmin = 1E-12
+ tnom = 30 ute = -1.379977 lute = 8.596947E-8
+ wute = 9.398486E-8 pute = -6.080689E-14 kt1 = -0.37073
+ kt1l = 0 kt2 = -0.019151 ua1 = 2.0117E-9
+ ub1 = -1.8012E-18 uc1 = -5.9821E-11 at = 5.302005E4
+ lat = -1.55406E-2 wat = -1.69896E-2 pat = 1.099201E-8
+ prt = 0 njs = 1.0773 xtis = 0.76
+ tpb = 1.344E-3 tpbsw = 9.9005E-4 tpbswg = 0
+ tcj = 6.7434E-4 tcjsw = 2.493E-4 tcjswg = 0
+ tvoff = 0 tvfbsdoff = 0 saref = 2.41E-6
+ sbref = 2.41E-6 wlod = 0 ku0 = -4.5E-8
+ kvsat = 0.3 kvth0 = 1.1E-8 tku0 = 0
+ llodku0 = 0 wlodku0 = 1 llodvth = 0
+ wlodvth = 1 lku0 = 0 wku0 = 2E-7
+ pku0 = 0 lkvth0 = 0 wkvth0 = 6.5E-7
+ pkvth0 = 0 stk2 = 0 lodk2 = 1
+ steta0 = 0 lodeta0 = 1

.model nhv_model.56 nmos
+ level = 54 lmin = 5E-7 lmax = 6E-7 wmin = 4.2E-7
+ wmax = 7.5E-7 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 1.16E-8
+ toxm = 1.16E-8 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 1E23 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {2.1346E-8+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {7.6507E-8-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = -4.1292E-9 dwb = -1.6944E-9 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = 0.790408 lvth0 = 1.726149E-8
+ wvth0 = 2.186923E-8 pvth0 = -1.465884E-14 k1 = 0.88325
+ k2 = -1.45094E-2 lk2 = -4.939263E-9 wk2 = 1.748426E-10
+ pk2 = 1.902463E-15 k3 = -0.884 k3b = 0.43
+ w0 = 0 lpe0 = 2.5E-8 lpeb = -2.182E-7
+ vbm = -3 dvtp0 = 0 dvtp1 = 0
+ dvt0 = 0 dvt1 = 0.53 dvt2 = -0.19251
+ dvt0w = 0.16 dvt1w = 6.9091E6 dvt2w = -0.036016
+ vfbsdoff = 0 u0 = 1.57162E-2 lu0 = 9.315056E-9
+ wu0 = 1.131059E-8 pu0 = -3.275241E-15 ua = -4.550441E-10
+ lua = 1.140487E-16 wua = 2.051982E-16 pua = -7.395696E-23
+ ub = -2.139209E-18 lub = 1.699652E-24 wub = 1.175569E-24
+ pub = -4.636969E-31 uc = 1.761389E-10 luc = -4.793193E-17
+ wuc = -2.802195E-17 puc = 9.723224E-24 ud = 0
+ up = 0 lp = 1 eu = 1.67
+ vsat = 7.734008E4 lvsat = 1.22221E-2 wvsat = 8.734194E-3
+ pvsat = -2.130279E-9 a0 = 1.1222 ags = 0.16025
+ b0 = 3.2933E-8 b1 = 0 keta = 4.85744E-2
+ lketa = -2.05535E-8 wketa = -2.23496E-8 pketa = 7.754998E-15
+ a1 = 0 a2 = 0.659726 rdsw = 724.62
+ rdswmin = 0 rdw = 0 rdwmin = 0
+ rsw = 0 rswmin = 0 prwb = 0.05626
+ prwg = 0.048 wr = 1 voff = -0.20613
+ voffl = -4.257949E-7 minv = 0 nfactor = 0.978922
+ lnfactor = 3.826528E-8 wnfactor = -7.503576E-8 pnfactor = 2.08086E-14
+ eta0 = 0.032 etab = -0.01932 dsub = 0.504
+ cit = -8E-4 cdsc = 0 cdscb = 0
+ cdscd = 0 pclm = -0.153668 lpclm = 3.258368E-7
+ wpclm = 4.486735E-7 ppclm = -3.311315E-14 pdiblc1 = 0.21098
+ pdiblc2 = 2E-4 pdiblcb = -0.26831 drout = 0.36075
+ pscbe1 = 9.3731E8 pscbe2 = 1.68E-6 pvag = 1.99
+ delta = 0.0246 fprout = 10.125 pdits = 0
+ pditsl = 0 pditsd = 0 lambda = 0
+ vtl = 0 lc = 5E-9 xn = 3
+ alpha0 = 2.089371E-4 lalpha0 = -6.747841E-11 walpha0 = -8.118268E-11
+ palpha0 = 2.816925E-17 alpha1 = 0 beta0 = 52.976772
+ lbeta0 = -5.557596E-6 wbeta0 = -1.132879E-5 pbeta0 = 3.930932E-12
+ aigbacc = 1 bigbacc = 0 cigbacc = 0
+ nigbacc = 1 aigbinv = 0.35 bigbinv = 0.03
+ cigbinv = 6E-3 eigbinv = 1.1 nigbinv = 3
+ aigc = 0.43 bigc = 0.054 cigc = 0.075
+ aigsd = 0.43 bigsd = 0.054 cigsd = 0.075
+ dlcig = 0 nigc = 1 poxedge = 1
+ pigcd = 1 ntox = 1 toxref = 1.16E-8
+ agidl = 5.06E-11 bgidl = 1.058E9 cgidl = 4E3
+ egidl = 0.8 noia = 2.6E41 noib = 0
+ noic = 0 em = 4.1E7 af = 1
+ ef = 0.89 kf = 0 lintnoi = 0
+ tnoia = 7.5E6 tnoib = 7.2E6 ntnoi = 1
+ rnoia = 0.794 rnoib = 0.38 xpart = 0
+ cgso = {2.754679E-10/sw_func_tox_hv_ratio} cgdo = {2.754679E-10/sw_func_tox_hv_ratio} cgbo = {0/sw_func_tox_hv_ratio}
+ ckappas = 0.6 cf = 0 clc = 1E-7
+ cle = 0.6 dlc = 6.5995E-8 dwc = 0
+ vfbcv = -1 noff = 4 voffcv = -0.4104
+ acde = 0.4176 moin = 15 cgsl = {4.49025E-11/sw_func_tox_hv_ratio}
+ cgdl = {4.49025E-11/sw_func_tox_hv_ratio} ijthsrev = 0.1 ijthsfwd = 0.1
+ xjbvs = 1 bvs = 12.636 jss = 3.75E-4
+ jsws = 5.84E-11 cjs = {8.310E-04*sw_func_nsd_pw_cj} mjs = 0.295
+ mjsws = 0.037586 cjsws = {8.643094E-11*sw_func_nsd_pw_cj} cjswgs = {5.47776E-11*sw_func_nsd_pw_cj}
+ mjswgs = 0.78692 pbs = 0.72468 pbsws = 0.29067
+ pbswgs = 0.54958 xrcrg1 = 12 xrcrg2 = 1
+ rbpb = 50 rbpd = 50 rbps = 50
+ rbdb = 50 rbsb = 50 gbmin = 1E-12
+ tnom = 30 ute = -1.961357 lute = 3.458381E-7
+ wute = 2.492201E-7 pute = -1.301949E-13 kt1 = -0.380618
+ lkt1 = 4.419726E-9 wkt1 = -4.209145E-8 pkt1 = 1.881429E-14
+ kt1l = 0 kt2 = -0.019151 ua1 = -1.43283E-9
+ lua1 = 1.539657E-15 ub1 = -8.069275E-18 lub1 = 2.801742E-24
+ wub1 = 4.919648E-24 pub1 = -2.199014E-30 uc1 = -5.9821E-11
+ at = -2.578625E4 lat = 1.96847E-2 wat = 9.554879E-3
+ pat = -8.729829E-10 prt = 0 njs = 1.0773
+ xtis = 0.76 tpb = 1.344E-3 tpbsw = 9.9005E-4
+ tpbswg = 0 tcj = 6.7434E-4 tcjsw = 2.493E-4
+ tcjswg = 0 tvoff = 0 tvfbsdoff = 0
+ saref = 2.02E-6 sbref = 2.01E-6 wlod = 0
+ ku0 = -4.5E-8 kvsat = 0.3 kvth0 = 1.1E-8
+ tku0 = 0 llodku0 = 0 wlodku0 = 1
+ llodvth = 0 wlodvth = 1 lku0 = 0
+ wku0 = 2E-7 pku0 = 0 lkvth0 = 0
+ wkvth0 = 6.5E-7 pkvth0 = 0 stk2 = 0
+ lodk2 = 1 steta0 = 0 lodeta0 = 1
.ends sky130_fd_pr__nfet_g5v0d10v5
