* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

******************************************************************
******************************************************************
*  *****************************************************
*  01/04/2022 Usman Suriono
*      Why     : Leakage corner was too low.
*      What    : Add variation to DIBL (deleta0) as the function of VT.
*  04/14/2021 Usman Suriono
*      Why     : New scalable sky130_fd_pr__nfet_01v8 model
*      What    : Converted from discrete nshort model
*                Replaced rsh from 1 to calculated rsh from the original model.
*                PDK netlist nrd/nrs = ratio of distance the middle of the contact to Gate.
*
*  *****************************************************
*
*  Nmos Model
*  -----------------------------------------------------

.subckt  sky130_fd_pr__nfet_01v8  d g s b  mult=1
+ 
.param  l = 1 w = 1 nf = 1 ad = 0 as = 0 pd = 0 ps = 0 nrd = {0.14/w} nrs = {0.14/w}
+ sa = 0 sb = 0 sd = 0
+ swx_vth = {sw_vth0_sky130_fd_pr__nfet_01v8+sw_mm_vth0_sky130_fd_pr__nfet_01v8*mismatch_factor*MC_MM_SWITCH*AGAUSS(0,1.0,1)/sqrt(l*w*mult)+sw_vth0_sky130_fd_pr__nfet_01v8_mc}
+ swx_nrds = {89.1*nf/w+443.5}

Msky130_fd_pr__nfet_01v8  d g s b nshort_model l = {l} w = {w} ad = {ad} as = {as} pd = {pd} ps = {ps} nrd = {nrd} nrs = {nrs} sa = {sa} sb = {sb} sd = {sd} nf = {nf}
* + deltox = 0.3*(sw_tox_lv_corner - sw_tox_lv_nom) + sw_tox_lv_mc + sw_mm_tox_lv * mismatch_factor*MC_MM_SWITCH*AGAUSS(0,1.0,1)/sqrt(l*w*mult)
* + mulu0  = sw_u0_sky130_fd_pr__nfet_01v8
+ delvto = {swx_vth*(0.008*8/l+0.992)*(0.035*7/w+0.965)*(0.001*56/(w*l)+0.999)}
* + mulvsat = sw_vsat_sky130_fd_pr__nfet_01v8
* + deleta0 = max(0,sw_vth0_sky130_fd_pr__nfet_01v8*2.8)



.model nshort_model.1 nmos
+ level = 54 lmin = 8E-6 lmax = 2.02E-5 wmin = 7E-6
+ wmax = 1.01E-3 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 4.148E-9
+ toxm = 4.148E-9 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 9.999999999999999E22 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {2.1859E-8+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {1.1932E-8-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = 0 dwb = 0 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = 0.5190093 k1 = 0.54086565
+ k2 = -0.026724591 k3 = 2 k3b = 0.54
+ w0 = 0 lpe0 = 1.0325E-7 lpeb = -7.082E-8
+ vbm = -3 dvtp0 = 0 dvtp1 = 0
+ dvt0 = 0 dvt1 = 0.53 dvt2 = -0.032
+ dvt0w = -3.58 dvt1w = 1.6706E6 dvt2w = 0.068
+ vfbsdoff = 0 u0 = 0.0318614 ua = -7.586635699999999E-10
+ ub = 1.674192E-18 uc = 4.9242E-11 ud = 0
+ up = 0 lp = 1 eu = 1.67
+ vsat = 8E4 a0 = 1.334619 ags = 0.4051693
+ b0 = 0 b1 = 2.1073424E-24 keta = -8.7946E-3
+ a1 = 0 a2 = 0.42385546 rdsw = 65.968
+ rdswmin = 0 rdw = 0 rdwmin = 0
+ rsw = 0 rswmin = 0 prwb = 0
+ prwg = 0.021507 wr = 1 voff = -0.1052686
+ voffl = 5.8197729E-9 minv = 0 nfactor = 2.63331
+ eta0 = 0.08 etab = -0.07 dsub = 0.56
+ cit = 0 cdsc = 0 cdscb = 0
+ cdscd = 5.4E-3 pclm = 0.026316 pdiblc1 = 0.39
+ pdiblc2 = 3.0734587E-3 pdiblcb = -0.025 drout = 0.56
+ pscbe1 = 7.5467416E8 pscbe2 = 1E-12 pvag = 0
+ delta = 0.01 fprout = 0 pdits = 0
+ pditsl = 0 pditsd = 0 lambda = 0
+ vtl = 0 lc = 5E-9 xn = 3
+ alpha0 = 3E-8 alpha1 = 0.85 beta0 = 13.86
+ aigbacc = 1 bigbacc = 0 cigbacc = 0
+ nigbacc = 0 aigbinv = 0.35 bigbinv = 0.03
+ cigbinv = 6E-3 eigbinv = 1.1 nigbinv = 0
+ aigc = 0.43 bigc = 0.054 cigc = 0.075
+ aigsd = 0.43 bigsd = 0.054 cigsd = 0.075
+ dlcig = 0 nigc = 0 poxedge = 1
+ pigcd = 1 ntox = 1 toxref = 4.148E-9
+ agidl = 0 bgidl = 2.3E9 cgidl = 0.5
+ egidl = 0.8 noia = 2.5E42 noib = 0
+ noic = 0 em = 4.1E7 af = 1
+ ef = 0.84 kf = 0 lintnoi = -1E-7
+ tnoia = 1.5E7 tnoib = 9.9E6 ntnoi = 1
+ rnoia = 0.94 rnoib = 0.26 xpart = 0
+ cgso = {2.449068E-10/sw_func_tox_lv_ratio} cgdo = {2.449068E-10/sw_func_tox_lv_ratio} cgbo = {1E-13/sw_func_tox_lv_ratio}
+ ckappas = 0.6 cf = 1.4067E-12 clc = 1E-7
+ cle = 0.6 dlc = 9.87908E-9 dwc = 0
+ vfbcv = -1 noff = 3.4037 voffcv = -0.17287
+ acde = 0.4 moin = 6.9 cgsl = {0/sw_func_tox_lv_ratio}
+ cgdl = {0/sw_func_tox_lv_ratio} ijthsrev = 0.1 ijthsfwd = 0.1
+ xjbvs = 1 bvs = 11.7 jss = 2.75E-3
+ jsws = 6E-10 cjs = {sw_nsd_pw_cj} mjs = 0.44
+ mjsws = 9E-4 cjsws = {3.67354204E-11*sw_func_nsd_pw_cj} cjswgs = {2.38232788E-10*sw_func_nsd_pw_cj}
+ mjswgs = 0.8 pbs = 0.729 pbsws = 0.2
+ pbswgs = 0.95578 xrcrg1 = 12 xrcrg2 = 1
+ rbpb = 50 rbpd = 50 rbps = 50
+ rbdb = 50 rbsb = 50 gbmin = 1E-12
+ tnom = 30 ute = -1.8134 kt1 = -0.31303
+ kt1l = 0 kt2 = -0.045313337 ua1 = 3.7602E-10
+ ub1 = -6.3962E-19 uc1 = 1.5829713E-11 at = 1.4E5
+ prt = 0 njs = 1.2928 xtis = 2
+ tpb = 1.2287E-3 tpbsw = 0 tpbswg = 0
+ tcj = 7.92E-4 tcjsw = 1E-5 tcjswg = 0
+ tvoff = 0 tvfbsdoff = 0 saref = 3E-6
+ sbref = 3E-6 wlod = 0 ku0 = -2.7E-8
+ kvsat = 0.2 kvth0 = 9.8E-9 tku0 = 0
+ llodku0 = 0 wlodku0 = 1 llodvth = 0
+ wlodvth = 1 lku0 = 0 wku0 = 0
+ pku0 = 0 lkvth0 = 0 wkvth0 = 2E-7
+ pkvth0 = 0 stk2 = 0 lodk2 = 1
+ steta0 = 0 lodeta0 = 1

.model nshort_model.2 nmos
+ level = 54 lmin = 4E-6 lmax = 8E-6 wmin = 7E-6
+ wmax = 1.01E-3 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 4.148E-9
+ toxm = 4.148E-9 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 9.999999999999999E22 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {2.1859E-8+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {1.1932E-8-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = 0 dwb = 0 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = 0.512816965197 lvth0 = 4.939090454626121E-8
+ k1 = 0.5317726245816 lk1 = 7.252720738861557E-8 k2 = -0.020817331231724
+ lk2 = -4.711710729909788E-8 k3 = 2 k3b = 0.54
+ w0 = 0 lpe0 = 1.0325E-7 lpeb = -7.082E-8
+ vbm = -3 dvtp0 = 0 dvtp1 = 0
+ dvt0 = 0 dvt1 = 0.53 dvt2 = -0.032
+ dvt0w = -3.58 dvt1w = 1.6706E6 dvt2w = 0.068
+ vfbsdoff = 0 u0 = 0.0321778010222 lu0 = -2.523657583606224E-9
+ ua = -7.638052605666998E-10 lua = 4.101082322991529E-17 ub = 1.702279424704E-18
+ lub = -2.240291193288636E-25 uc = 5.555113379800001E-11 luc = -5.032250921504456E-17
+ ud = 0 up = 0 lp = 1
+ eu = 1.67 vsat = 8E4 a0 = 1.42994189043
+ la0 = -7.603083379827791E-7 ags = 0.3924181300582 lags = 1.017050656149089E-7
+ b0 = 0 b1 = 4.202112395241601E-24 lb1 = -1.670817037076636E-29
+ keta = -0.0155666554318 lketa = 5.401483512357553E-8 a1 = 0
+ a2 = 0.42385546 rdsw = 65.968 rdswmin = 0
+ rdw = 0 rdwmin = 0 rsw = 0
+ rswmin = 0 prwb = 0 prwg = 0.021507
+ wr = 1 voff = -0.10886654582436 lvoff = 2.869770521572751E-8
+ voffl = 5.8197729E-9 minv = 0 nfactor = 2.59233591852
+ lnfactor = 3.268148463595616E-7 eta0 = 0.08 etab = -0.07
+ dsub = 0.56 cit = 0 cdsc = 0
+ cdscb = 0 cdscd = 5.4E-3 pclm = -0.531042839936
+ lpclm = 4.445569908131768E-6 pdiblc1 = 0.39 pdiblc2 = 3.0564335814718E-3
+ lpdiblc2 = 1.357946607970441E-10 pdiblcb = -0.025 drout = 0.56
+ pscbe1 = 7.0961873396144E8 lpscbe1 = 359.36820562149586 pscbe2 = 1E-12
+ pvag = 0 delta = 0.01 fprout = 0
+ pdits = 0 pditsl = 0 pditsd = 0
+ lambda = 0 vtl = 0 lc = 5E-9
+ xn = 3 alpha0 = 3E-8 alpha1 = 0.85
+ beta0 = 13.86 aigbacc = 1 bigbacc = 0
+ cigbacc = 0 nigbacc = 0 aigbinv = 0.35
+ bigbinv = 0.03 cigbinv = 6E-3 eigbinv = 1.1
+ nigbinv = 0 aigc = 0.43 bigc = 0.054
+ cigc = 0.075 aigsd = 0.43 bigsd = 0.054
+ cigsd = 0.075 dlcig = 0 nigc = 0
+ poxedge = 1 pigcd = 1 ntox = 1
+ toxref = 4.148E-9 agidl = 0 bgidl = 2.3E9
+ cgidl = 0.5 egidl = 0.8 noia = 2.5E42
+ noib = 0 noic = 0 em = 4.1E7
+ af = 1 ef = 0.84 kf = 0
+ lintnoi = -1E-7 tnoia = 1.5E7 tnoib = 9.9E6
+ ntnoi = 1 rnoia = 0.94 rnoib = 0.26
+ xpart = 0 cgso = {2.449068E-10/sw_func_tox_lv_ratio} cgdo = {2.449068E-10/sw_func_tox_lv_ratio}
+ cgbo = {1E-13/sw_func_tox_lv_ratio} ckappas = 0.6 cf = 1.4067E-12
+ clc = 1E-7 cle = 0.6 dlc = 9.87908E-9
+ dwc = 0 vfbcv = -1 noff = 3.4037
+ voffcv = -0.17287 acde = 0.4 moin = 6.9
+ cgsl = {0/sw_func_tox_lv_ratio} cgdl = {0/sw_func_tox_lv_ratio} ijthsrev = 0.1
+ ijthsfwd = 0.1 xjbvs = 1 bvs = 11.7
+ jss = 2.75E-3 jsws = 6E-10 cjs = {sw_nsd_pw_cj}
+ mjs = 0.44 mjsws = 9E-4 cjsws = {3.67354204E-11*sw_func_nsd_pw_cj}
+ cjswgs = {2.38232788E-10*sw_func_nsd_pw_cj} mjswgs = 0.8 pbs = 0.729
+ pbsws = 0.2 pbswgs = 0.95578 xrcrg1 = 12
+ xrcrg2 = 1 rbpb = 50 rbpd = 50
+ rbps = 50 rbdb = 50 rbsb = 50
+ gbmin = 1E-12 tnom = 30 ute = -1.7738374468
+ lute = -3.155563048304357E-7 kt1 = -0.31093258826 lkt1 = -1.672924128623665E-8
+ kt1l = 0 kt2 = -0.04419860739172 lkt2 = -8.891234958867991E-9
+ ua1 = 5.718049366400001E-10 lua1 = -1.561607281392023E-15 ub1 = -8.959316669E-19
+ lub1 = 2.044376713581099E-24 uc1 = 1.388679293995998E-12 luc1 = 1.151836488196719E-16
+ at = 1.4E5 prt = 0 njs = 1.2928
+ xtis = 2 tpb = 1.2287E-3 tpbsw = 0
+ tpbswg = 0 tcj = 7.92E-4 tcjsw = 1E-5
+ tcjswg = 0 tvoff = 0 tvfbsdoff = 0
+ saref = 3E-6 sbref = 3E-6 wlod = 0
+ ku0 = -2.7E-8 kvsat = 0.2 kvth0 = 9.8E-9
+ tku0 = 0 llodku0 = 0 wlodku0 = 1
+ llodvth = 0 wlodvth = 1 lku0 = 0
+ wku0 = 0 pku0 = 0 lkvth0 = 0
+ wkvth0 = 2E-7 pkvth0 = 0 stk2 = 0
+ lodk2 = 1 steta0 = 0 lodeta0 = 1

.model nshort_model.3 nmos
+ level = 54 lmin = 2E-6 lmax = 4E-6 wmin = 7E-6
+ wmax = 1.01E-3 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 4.148E-9
+ toxm = 4.148E-9 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 9.999999999999999E22 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {2.1859E-8+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {1.1932E-8-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = 0 dwb = 0 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = 0.518547603504 lvth0 = 2.660510727081945E-8
+ k1 = 0.55001325 k2 = -0.031298059138892 lk2 = -5.444307761202527E-9
+ k3 = 2 k3b = 0.54 w0 = 0
+ lpe0 = 1.0325E-7 lpeb = -7.082E-8 vbm = -3
+ dvtp0 = 0 dvtp1 = 0 dvt0 = 0
+ dvt1 = 0.53 dvt2 = -0.032 dvt0w = -3.58
+ dvt1w = 1.6706E6 dvt2w = 0.068 vfbsdoff = 0
+ u0 = 0.0332068088984 lu0 = -6.615132844448578E-9 ua = -5.832601931146001E-10
+ lua = -6.768609190888065E-16 ub = 1.523794986112E-18 lub = 4.856492823965773E-25
+ uc = 1.185089150800001E-11 luc = 1.234355973629469E-16 ud = 0
+ up = 0 lp = 1 eu = 1.67
+ vsat = 8E4 a0 = 1.249866442836 la0 = -4.430386808816161E-8
+ ags = 0.254250418768 lags = 6.510786765134796E-7 b0 = 0
+ b1 = 0 keta = -3.814351151439999E-3 lketa = 7.286074991482034E-9
+ a1 = 0 a2 = 0.42385546 rdsw = 65.968
+ rdswmin = 0 rdw = 0 rdwmin = 0
+ rsw = 0 rswmin = 0 prwb = 0
+ prwg = 0.021507 wr = 1 voff = -0.10138368469656
+ lvoff = -1.055168297518725E-9 voffl = 5.8197729E-9 minv = 0
+ nfactor = 2.59433840112 lnfactor = 3.188527032043281E-7 eta0 = 0.158551406
+ leta0 = -3.123310732472159E-7 etab = -0.138670043175847 letab = 2.730414307930405E-7
+ dsub = 0.8564204 ldsub = -1.1786078235744E-6 cit = 0
+ cdsc = 0 cdscb = 0 cdscd = 5.4E-3
+ pclm = 0.61455745516 lpclm = -1.094926668100615E-7 pdiblc1 = 0.39
+ pdiblc2 = 1.389224399096801E-3 lpdiblc2 = 6.764845110368845E-9 pdiblcb = -0.025
+ drout = 0.56 pscbe1 = 8E8 pscbe2 = 1E-12
+ pvag = 0 delta = 0.01 fprout = 0
+ pdits = 0 pditsl = 0 pditsd = 0
+ lambda = 0 vtl = 0 lc = 5E-9
+ xn = 3 alpha0 = 3E-8 alpha1 = 0.85
+ beta0 = 13.86 aigbacc = 1 bigbacc = 0
+ cigbacc = 0 nigbacc = 0 aigbinv = 0.35
+ bigbinv = 0.03 cigbinv = 6E-3 eigbinv = 1.1
+ nigbinv = 0 aigc = 0.43 bigc = 0.054
+ cigc = 0.075 aigsd = 0.43 bigsd = 0.054
+ cigsd = 0.075 dlcig = 0 nigc = 0
+ poxedge = 1 pigcd = 1 ntox = 1
+ toxref = 4.148E-9 agidl = 0 bgidl = 2.3E9
+ cgidl = 0.5 egidl = 0.8 noia = 2.5E42
+ noib = 0 noic = 0 em = 4.1E7
+ af = 1 ef = 0.84 kf = 0
+ lintnoi = -1E-7 tnoia = 1.5E7 tnoib = 9.9E6
+ ntnoi = 1 rnoia = 0.94 rnoib = 0.26
+ xpart = 0 cgso = {2.449068E-10/sw_func_tox_lv_ratio} cgdo = {2.449068E-10/sw_func_tox_lv_ratio}
+ cgbo = {1E-13/sw_func_tox_lv_ratio} ckappas = 0.6 cf = 1.4067E-12
+ clc = 1E-7 cle = 0.6 dlc = 9.87908E-9
+ dwc = 0 vfbcv = -1 noff = 3.4037
+ voffcv = -0.17287 acde = 0.4 moin = 6.9
+ cgsl = {0/sw_func_tox_lv_ratio} cgdl = {0/sw_func_tox_lv_ratio} ijthsrev = 0.1
+ ijthsfwd = 0.1 xjbvs = 1 bvs = 11.7
+ jss = 2.75E-3 jsws = 6E-10 cjs = {sw_nsd_pw_cj}
+ mjs = 0.44 mjsws = 9E-4 cjsws = {3.67354204E-11*sw_func_nsd_pw_cj}
+ cjswgs = {2.38232788E-10*sw_func_nsd_pw_cj} mjswgs = 0.8 pbs = 0.729
+ pbsws = 0.2 pbswgs = 0.95578 xrcrg1 = 12
+ xrcrg2 = 1 rbpb = 50 rbpd = 50
+ rbps = 50 rbdb = 50 rbsb = 50
+ gbmin = 1E-12 tnom = 30 ute = -1.9898498044
+ lute = 5.433382066677978E-7 kt1 = -0.30640547888 lkt1 = -3.472964386799237E-8
+ kt1l = 0 kt2 = -0.046434757 ua1 = -1.235654670399999E-10
+ lua1 = 1.203280014014557E-15 ub1 = -2.004199992800001E-19 lub1 = -7.210722664628177E-25
+ uc1 = 2.435133106997601E-11 luc1 = 2.388102243773389E-17 at = 1.6476098408E5
+ lat = -0.098453040195915 prt = 0 njs = 1.2928
+ xtis = 2 tpb = 1.2287E-3 tpbsw = 0
+ tpbswg = 0 tcj = 7.92E-4 tcjsw = 1E-5
+ tcjswg = 0 tvoff = 0 tvfbsdoff = 0
+ saref = 3E-6 sbref = 3E-6 wlod = 0
+ ku0 = -2.7E-8 kvsat = 0.2 kvth0 = 9.8E-9
+ tku0 = 0 llodku0 = 0 wlodku0 = 1
+ llodvth = 0 wlodvth = 1 lku0 = 0
+ wku0 = 0 pku0 = 0 lkvth0 = 0
+ wkvth0 = 2E-7 pkvth0 = 0 stk2 = 0
+ lodk2 = 1 steta0 = 0 lodeta0 = 1

.model nshort_model.4 nmos
+ level = 54 lmin = 1E-6 lmax = 2E-6 wmin = 7E-6
+ wmax = 1.01E-3 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 4.148E-9
+ toxm = 4.148E-9 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 9.999999999999999E22 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {2.1859E-8+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {1.1932E-8-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = 0 dwb = 0 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = 0.5080903920928 lvth0 = 4.72699792001026E-8
+ k1 = 0.51693995598888 lk1 = 6.510428271915861E-8 k2 = -0.021137344468272
+ lk2 = -2.552326180754284E-8 k3 = 2 k3b = 0.54
+ w0 = 0 lpe0 = 1.0325E-7 lpeb = -7.082E-8
+ vbm = -3 dvtp0 = 0 dvtp1 = 0
+ dvt0 = 0 dvt1 = 0.53 dvt2 = -0.032
+ dvt0w = -3.58 dvt1w = 1.6706E6 dvt2w = 0.068
+ vfbsdoff = 0 u0 = 0.0337134753824 lu0 = -7.616374723474404E-9
+ ua = -4.202807300495199E-10 lua = -9.98930503312382E-16 ub = 1.303723306488E-18
+ lub = 9.205408510820295E-25 uc = 8.743424397599998E-11 luc = -2.592738644975672E-17
+ ud = 0 up = 0 lp = 1
+ eu = 1.67 vsat = 6.018443919999999E4 lvsat = 0.039158243057069
+ a0 = 1.365388682704 la0 = -2.725915250919517E-7 ags = 0.281209620648
+ lags = 5.978036271471438E-7 b0 = 0 b1 = 0
+ keta = 0.063267337619048 lketa = -1.252764651286751E-7 a1 = 0
+ a2 = 0.42385546 rdsw = 65.968 rdswmin = 0
+ rdw = 0 rdwmin = 0 rsw = 0
+ rswmin = 0 prwb = 0 prwg = 0.021507
+ wr = 1 voff = -0.08364582852264 lvoff = -3.610758444562427E-8
+ voffl = 5.8197729E-9 minv = 0 nfactor = 2.8687414836808
+ lnfactor = -2.234051067550413E-7 eta0 = -1.482776250000001E-3 leta0 = 3.918235527570001E-9
+ etab = -6.8439114830552E-4 letab = 3.630163379423571E-10 dsub = 0.26
+ cit = 0 cdsc = 0 cdscb = 0
+ cdscd = 5.4E-3 pclm = 0.72262349592 lpclm = -3.230458603333653E-7
+ pdiblc1 = 0.0804062659 lpdiblc1 = 6.117993233294377E-7 pdiblc2 = 5.594452912790401E-3
+ lpdiblc2 = -1.545258343767571E-9 pdiblcb = -0.049216379985545 lpdiblcb = 4.785486027911472E-8
+ drout = 0.8528408 ldrout = -5.786932471488001E-7 pscbe1 = 1.32606452329984E9
+ lpscbe1 = -1.039575042815653E3 pscbe2 = 1E-12 pvag = 0
+ delta = 0.01 fprout = 0 pdits = 0
+ pditsl = 0 pditsd = 0 lambda = 0
+ vtl = 0 lc = 5E-9 xn = 3
+ alpha0 = -2.51771496E-6 lalpha0 = 5.03463125019456E-12 alpha1 = 0.816811376
+ lalpha1 = 6.558523467686407E-8 beta0 = 11.154151007999996 lbeta0 = 5.347125603654916E-6
+ aigbacc = 1 bigbacc = 0 cigbacc = 0
+ nigbacc = 0 aigbinv = 0.35 bigbinv = 0.03
+ cigbinv = 6E-3 eigbinv = 1.1 nigbinv = 0
+ aigc = 0.43 bigc = 0.054 cigc = 0.075
+ aigsd = 0.43 bigsd = 0.054 cigsd = 0.075
+ dlcig = 0 nigc = 0 poxedge = 1
+ pigcd = 1 ntox = 1 toxref = 4.148E-9
+ agidl = 0 bgidl = 2.3E9 cgidl = 0.5
+ egidl = 0.8 noia = 2.5E42 noib = 0
+ noic = 0 em = 4.1E7 af = 1
+ ef = 0.84 kf = 0 lintnoi = -1E-7
+ tnoia = 1.5E7 tnoib = 9.9E6 ntnoi = 1
+ rnoia = 0.94 rnoib = 0.26 xpart = 0
+ cgso = {2.449068E-10/sw_func_tox_lv_ratio} cgdo = {2.449068E-10/sw_func_tox_lv_ratio} cgbo = {1E-13/sw_func_tox_lv_ratio}
+ ckappas = 0.6 cf = 1.4067E-12 clc = 1E-7
+ cle = 0.6 dlc = 9.87908E-9 dwc = 0
+ vfbcv = -1 noff = 3.4037 voffcv = -0.17287
+ acde = 0.4 moin = 6.9 cgsl = {0/sw_func_tox_lv_ratio}
+ cgdl = {0/sw_func_tox_lv_ratio} ijthsrev = 0.1 ijthsfwd = 0.1
+ xjbvs = 1 bvs = 11.7 jss = 2.75E-3
+ jsws = 6E-10 cjs = {sw_nsd_pw_cj} mjs = 0.44
+ mjsws = 9E-4 cjsws = {3.67354204E-11*sw_func_nsd_pw_cj} cjswgs = {2.38232788E-10*sw_func_nsd_pw_cj}
+ mjswgs = 0.8 pbs = 0.729 pbsws = 0.2
+ pbswgs = 0.95578 xrcrg1 = 12 xrcrg2 = 1
+ rbpb = 50 rbpd = 50 rbps = 50
+ rbdb = 50 rbsb = 50 gbmin = 1E-12
+ tnom = 30 ute = -2.52321946026608 lute = 1.59734918493237E-6
+ kt1 = -0.37404601544 lkt1 = 9.893725548753985E-8 kt1l = 0
+ kt2 = -0.066031623371848 lkt2 = 3.869874711599023E-8 ua1 = -1.1925068841624E-9
+ lua1 = 3.315653630281149E-15 ub1 = 3.155993453608003E-19 lub1 = -1.74079667010391E-24
+ uc1 = 1.7468532419304E-11 luc1 = 3.748236863207827E-17 at = 1.65283238064E5
+ lat = -0.099485085094841 prt = 0 njs = 1.2928
+ xtis = 2 tpb = 1.2287E-3 tpbsw = 0
+ tpbswg = 0 tcj = 7.92E-4 tcjsw = 1E-5
+ tcjswg = 0 tvoff = 0 tvfbsdoff = 0
+ saref = 3E-6 sbref = 3E-6 wlod = 0
+ ku0 = -2.7E-8 kvsat = 0.2 kvth0 = 9.8E-9
+ tku0 = 0 llodku0 = 0 wlodku0 = 1
+ llodvth = 0 wlodvth = 1 lku0 = 0
+ wku0 = 0 pku0 = 0 lkvth0 = 0
+ wkvth0 = 2E-7 pkvth0 = 0 stk2 = 0
+ lodk2 = 1 steta0 = 0 lodeta0 = 1

.model nshort_model.5 nmos
+ level = 54 lmin = 5E-7 lmax = 1E-6 wmin = 7E-6
+ wmax = 1.01E-3 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 4.148E-9
+ toxm = 4.148E-9 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 9.999999999999999E22 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {2.1859E-8+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {1.1932E-8-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = 0 dwb = 0 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = 0.5382094278448 lvth0 = 1.786970411728827E-8
+ k1 = 0.67685538541968 lk1 = -9.099492490370467E-8 k2 = -0.084108743215152
+ lk2 = 3.59453874796416E-8 k3 = 2 k3b = 0.54
+ w0 = 0 lpe0 = 1.0325E-7 lpeb = -7.082E-8
+ vbm = -3 dvtp0 = 0 dvtp1 = 0
+ dvt0 = 0 dvt1 = 0.53 dvt2 = -0.032
+ dvt0w = -3.58 dvt1w = 1.6706E6 dvt2w = 0.068
+ vfbsdoff = 0 u0 = 0.028060177904 lu0 = -2.097987536098945E-9
+ ua = -1.287815499504323E-9 lua = -1.520985835958479E-16 ub = 2.22680937888E-18
+ lub = 1.948330472159232E-26 uc = 4.004109772800001E-11 luc = 2.033476975618098E-17
+ ud = 0 up = 0 lp = 1
+ eu = 1.67 vsat = 8.75341272496E4 lvsat = 0.012461227963084
+ a0 = 0.692019044176 la0 = 3.84708820382216E-7 ags = 0.554264922816
+ lags = 3.31264516710081E-7 b0 = 0 b1 = 0
+ keta = -0.101468423037136 lketa = 3.552804133520978E-8 a1 = 0
+ a2 = 0.42385546 rdsw = 65.968 rdswmin = 0
+ rdw = 0 rdwmin = 0 rsw = 0
+ rswmin = 0 prwb = 0 prwg = 0.021507
+ wr = 1 voff = -0.10764602671632 lvoff = -1.268012698163826E-8
+ voffl = 5.8197729E-9 minv = 0 nfactor = 2.4855724494352
+ lnfactor = 1.506199816573214E-7 eta0 = -0.4616715915 leta0 = 4.531251048904439E-7
+ etab = -3.125E-4 dsub = 0.13096570606928 ldsub = 1.259550195403573E-7
+ cit = 0 cdsc = 0 cdscb = 0
+ cdscd = 5.4E-3 pclm = 0.25367674176 lpclm = 1.347099484853606E-7
+ pdiblc1 = 0.4283015482 lpdiblc1 = 2.722062140462447E-7 pdiblc2 = 4.5695576175984E-3
+ lpdiblc2 = -5.448211499000314E-10 pdiblcb = 0.02343275997109 lpdiblcb = -2.306058060159479E-8
+ drout = 0.03264278406992 ldrout = 2.219315633291245E-7 pscbe1 = -2.436478200319994E7
+ lpscbe1 = 278.6276175456356 pscbe2 = 1E-12 pvag = 0
+ delta = 0.01 fprout = 0 pdits = 0
+ pditsl = 0 pditsd = 0 lambda = 0
+ vtl = 0 lc = 5E-9 xn = 3
+ alpha0 = -5.596339199999991E-7 lalpha0 = 3.123277856133119E-12 alpha1 = 0.916377248
+ lalpha1 = -3.160459735372802E-8 beta0 = 14.567474304000003 lbeta0 = 2.015257854790655E-6
+ aigbacc = 1 bigbacc = 0 cigbacc = 0
+ nigbacc = 0 aigbinv = 0.35 bigbinv = 0.03
+ cigbinv = 6E-3 eigbinv = 1.1 nigbinv = 0
+ aigc = 0.43 bigc = 0.054 cigc = 0.075
+ aigsd = 0.43 bigsd = 0.054 cigsd = 0.075
+ dlcig = 0 nigc = 0 poxedge = 1
+ pigcd = 1 ntox = 1 toxref = 4.148E-9
+ agidl = 0 bgidl = 2.3E9 cgidl = 0.5
+ egidl = 0.8 noia = 2.5E42 noib = 0
+ noic = 0 em = 4.1E7 af = 1
+ ef = 0.84 kf = 0 lintnoi = -1E-7
+ tnoia = 1.5E7 tnoib = 9.9E6 ntnoi = 1
+ rnoia = 0.94 rnoib = 0.26 xpart = 0
+ cgso = {2.449068E-10/sw_func_tox_lv_ratio} cgdo = {2.449068E-10/sw_func_tox_lv_ratio} cgbo = {1E-13/sw_func_tox_lv_ratio}
+ ckappas = 0.6 cf = 1.4067E-12 clc = 1E-7
+ cle = 0.6 dlc = 9.87908E-9 dwc = 0
+ vfbcv = -1 noff = 3.4037 voffcv = -0.17287
+ acde = 0.4 moin = 6.9 cgsl = {0/sw_func_tox_lv_ratio}
+ cgdl = {0/sw_func_tox_lv_ratio} ijthsrev = 0.1 ijthsfwd = 0.1
+ xjbvs = 1 bvs = 11.7 jss = 2.75E-3
+ jsws = 6E-10 cjs = {sw_nsd_pw_cj} mjs = 0.44
+ mjsws = 9E-4 cjsws = {3.67354204E-11*sw_func_nsd_pw_cj} cjswgs = {2.38232788E-10*sw_func_nsd_pw_cj}
+ mjswgs = 0.8 pbs = 0.729 pbsws = 0.2
+ pbswgs = 0.95578 xrcrg1 = 12 xrcrg2 = 1
+ rbpb = 50 rbpd = 50 rbps = 50
+ rbdb = 50 rbsb = 50 gbmin = 1E-12
+ tnom = 30 ute = -0.37232496106784 lute = -5.022163679370029E-7
+ kt1 = -0.26882377568 lkt1 = -3.773960742827527E-9 kt1l = 0
+ kt2 = -0.017158188825376 lkt2 = -9.008371788464771E-9 ua1 = 3.2341434902304E-9
+ lua1 = -1.005359159577142E-15 ub1 = -1.7234129065664E-18 lub1 = 2.495565934432993E-25
+ uc1 = 1.22134998482928E-10 luc1 = -6.468633688540339E-17 at = 7.282967913599999E4
+ lat = -9.237837897098495E-3 prt = 0 njs = 1.2928
+ xtis = 2 tpb = 1.2287E-3 tpbsw = 0
+ tpbswg = 0 tcj = 7.92E-4 tcjsw = 1E-5
+ tcjswg = 0 tvoff = 0 tvfbsdoff = 0
+ saref = 2.75E-6 sbref = 2.74E-6 wlod = 0
+ ku0 = -2.7E-8 kvsat = 0.2 kvth0 = 9.8E-9
+ tku0 = 0 llodku0 = 0 wlodku0 = 1
+ llodvth = 0 wlodvth = 1 lku0 = 0
+ wku0 = 0 pku0 = 0 lkvth0 = 0
+ wkvth0 = 2E-7 pkvth0 = 0 stk2 = 0
+ lodk2 = 1 steta0 = 0 lodeta0 = 1

.model nshort_model.6 nmos
+ level = 54 lmin = 2.5E-7 lmax = 5E-7 wmin = 7E-6
+ wmax = 1.01E-3 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 4.148E-9
+ toxm = 4.148E-9 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 9.999999999999999E22 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {2.1859E-8+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {1.1932E-8-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = 0 dwb = 0 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = 0.619842499536 lvth0 = -2.099874010547288E-8
+ k1 = 0.23608175037696 lk1 = 1.188732705909957E-7 k2 = 0.062088194974752
+ lk2 = -3.366423788234651E-8 k3 = 2 k3b = 0.54
+ w0 = 0 lpe0 = 1.0325E-7 lpeb = -7.082E-8
+ vbm = -3 dvtp0 = 0 dvtp1 = 0
+ dvt0 = 0 dvt1 = 0.53 dvt2 = -0.032
+ dvt0w = -3.58 dvt1w = 1.6706E6 dvt2w = 0.068
+ vfbsdoff = 0 u0 = 0.0291195166656 lu0 = -2.602376856692121E-9
+ ua = -1.131158186856954E-9 lua = -2.26688769810516E-16 ub = 1.96890384416E-18
+ lub = 1.422814144010342E-25 uc = 8.1085543584E-11 luc = 7.920314840885738E-19
+ ud = 0 up = 0 lp = 1
+ eu = 1.67 vsat = 9.20231471392E4 lvsat = 0.01032384398893
+ a0 = 1.5 ags = 2.363013351136 lags = -5.299457249564905E-7
+ b0 = 0 b1 = 0 keta = -0.016261925814048
+ lketa = -5.04183942660244E-9 a1 = 0 a2 = 0.42385546
+ rdsw = 65.968 rdswmin = 0 rdw = 0
+ rdwmin = 0 rsw = 0 rswmin = 0
+ prwb = 0 prwg = 0.021507 wr = 1
+ voff = -0.12699208835136 lvoff = -3.468770578976856E-9 voffl = 5.8197729E-9
+ minv = 0 nfactor = 2.781656050751999 lnfactor = 9.643920060745905E-9
+ eta0 = 0.49 etab = 2.097234539241599E-4 letab = -2.486493864576338E-10
+ dsub = 0.24857689844288 ldsub = 6.99560968483609E-8 cit = 0
+ cdsc = 0 cdscb = 0 cdscd = 5.4E-3
+ pclm = 0.64931522784 lpclm = -5.366777772282621E-8 pdiblc1 = 1.79766578554656
+ lpdiblc1 = -3.797973964669969E-7 pdiblc2 = 4.2262572879392E-3 lpdiblc2 = -3.813635041374189E-10
+ pdiblcb = 0.1559088 lpdiblcb = -8.61371923968E-8 drout = 0.04535187186016
+ ldrout = 2.158803091050309E-7 pscbe1 = 3.4447147080704E8 lpscbe1 = 103.0113994775792
+ pscbe2 = 1E-12 pvag = 0 delta = 0.01
+ fprout = 0 pdits = 0 pditsl = 0
+ pditsd = 0 lambda = 0 vtl = 0
+ lc = 5E-9 xn = 3 alpha0 = 9.03926784E-6
+ lalpha0 = -1.44710483226624E-12 alpha1 = 0.85 beta0 = 18.504214112000003
+ lbeta0 = 1.408343095687672E-7 aigbacc = 1 bigbacc = 0
+ cigbacc = 0 nigbacc = 0 aigbinv = 0.35
+ bigbinv = 0.03 cigbinv = 6E-3 eigbinv = 1.1
+ nigbinv = 0 aigc = 0.43 bigc = 0.054
+ cigc = 0.075 aigsd = 0.43 bigsd = 0.054
+ cigsd = 0.075 dlcig = 0 nigc = 0
+ poxedge = 1 pigcd = 1 ntox = 1
+ toxref = 4.148E-9 agidl = 0 bgidl = 2.3E9
+ cgidl = 0.5 egidl = 0.8 noia = 2.5E42
+ noib = 0 noic = 0 em = 4.1E7
+ af = 1 ef = 0.84 kf = 0
+ lintnoi = -1E-7 tnoia = 1.5E7 tnoib = 9.9E6
+ ntnoi = 1 rnoia = 0.94 rnoib = 0.26
+ xpart = 0 cgso = {2.449068E-10/sw_func_tox_lv_ratio} cgdo = {2.449068E-10/sw_func_tox_lv_ratio}
+ cgbo = {1E-13/sw_func_tox_lv_ratio} ckappas = 0.6 cf = 1.4067E-12
+ clc = 1E-7 cle = 0.6 dlc = 9.87908E-9
+ dwc = 0 vfbcv = -1 noff = 3.4037
+ voffcv = -0.17287 acde = 0.4 moin = 6.9
+ cgsl = {0/sw_func_tox_lv_ratio} cgdl = {0/sw_func_tox_lv_ratio} ijthsrev = 0.1
+ ijthsfwd = 0.1 xjbvs = 1 bvs = 11.7
+ jss = 2.75E-3 jsws = 6E-10 cjs = {sw_nsd_pw_cj}
+ mjs = 0.44 mjsws = 9E-4 cjsws = {3.67354204E-11*sw_func_nsd_pw_cj}
+ cjswgs = {2.38232788E-10*sw_func_nsd_pw_cj} mjswgs = 0.8 pbs = 0.729
+ pbsws = 0.2 pbswgs = 0.95578 xrcrg1 = 12
+ xrcrg2 = 1 rbpb = 50 rbpd = 50
+ rbps = 50 rbdb = 50 rbsb = 50
+ gbmin = 1E-12 tnom = 30 ute = -1.93202640173856
+ lute = 2.40413637218191E-7 kt1 = -0.26326140369024 lkt1 = -6.422406292543893E-9
+ kt1l = 0 kt2 = -0.032574405333824 lkt2 = -1.668156124998376E-9
+ ua1 = 8.170587259455999E-10 lua1 = 1.455019117503658E-16 ub1 = -1.5900272984864E-18
+ lub1 = 1.860469035545205E-25 uc1 = -1.0760097217472E-10 luc1 = 4.469922923964648E-17
+ at = 7.8306200981152E4 lat = -0.011845407102362 prt = 0
+ njs = 1.2928 xtis = 2 tpb = 1.2287E-3
+ tpbsw = 0 tpbswg = 0 tcj = 7.92E-4
+ tcjsw = 1E-5 tcjswg = 0 tvoff = 0
+ tvfbsdoff = 0 saref = 1.75E-6 sbref = 1.74E-6
+ wlod = 0 ku0 = -2.7E-8 kvsat = 0.2
+ kvth0 = 9.8E-9 tku0 = 0 llodku0 = 0
+ wlodku0 = 1 llodvth = 0 wlodvth = 1
+ lku0 = 0 wku0 = 0 pku0 = 0
+ lkvth0 = 0 wkvth0 = 2E-7 pkvth0 = 0
+ stk2 = 0 lodk2 = 1 steta0 = 0
+ lodeta0 = 1

.model nshort_model.7 nmos
+ level = 54 lmin = 1.8E-7 lmax = 2.5E-7 wmin = 7E-6
+ wmax = 1.01E-3 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 4.148E-9
+ toxm = 4.148E-9 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 9.999999999999999E22 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {2.1859E-8+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {1.1932E-8-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = 0 dwb = 0 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = 0.65652651648 lvth0 = -2.929431696112129E-8
+ k1 = 0.482996222366857 lk1 = 6.30370195530884E-8 k2 = -5.405528737371407E-3
+ lk2 = -1.840147717698178E-8 k3 = 2 k3b = 0.54
+ w0 = 0 lpe0 = 1.0325E-7 lpeb = -7.082E-8
+ vbm = -3 dvtp0 = 0 dvtp1 = 0
+ dvt0 = 0 dvt1 = 0.53 dvt2 = -0.032
+ dvt0w = -3.58 dvt1w = 1.6706E6 dvt2w = 0.068
+ vfbsdoff = 0 u0 = -9.249914388571437E-3 lu0 = 6.07433280417399E-9
+ ua = -5.182469379794288E-9 lua = 6.894585381155608E-16 ub = 4.782295578628572E-18
+ lub = -4.939277388647507E-25 uc = 8.054853862857142E-11 luc = 9.134676366893717E-19
+ ud = 0 up = 0 lp = 1
+ eu = 1.67 vsat = 1.143149747977143E5 lvsat = 5.282859249544082E-3
+ a0 = 1.5 ags = -2.725047682628572 lags = 6.206480449748947E-7
+ b0 = 0 b1 = 0 keta = -0.037026358549829
+ lketa = -3.462536654639678E-10 a1 = 0 a2 = 0.42385546
+ rdsw = 65.968 rdswmin = 0 rdw = 0
+ rdwmin = 0 rsw = 0 rswmin = 0
+ prwb = 0 prwg = 0.021507 wr = 1
+ voff = -0.11438617872 lvoff = -6.319420559374082E-9 voffl = 5.8197729E-9
+ minv = 0 nfactor = 2.064372182194286 lnfactor = 1.718476249609129E-7
+ eta0 = 1.513844491134514 leta0 = -2.315280978471945E-7 etab = 0.060377227297585
+ letab = -1.385468803564775E-8 dsub = 0.912559318723429 ldsub = -8.019423174420126E-8
+ cit = 0 cdsc = 0 cdscb = 0
+ cdscd = 8.522720000000001E-3 lcdscd = -7.061594099200002E-10 pclm = 0.692053373714286
+ lpclm = -6.333241107825373E-8 pdiblc1 = -0.454454416598857 lpdiblc1 = 1.294880575653592E-7
+ pdiblc2 = -0.011489398761726 lpdiblc2 = 3.172512092309606E-9 pdiblcb = -0.534247159427886
+ lpdiblcb = 6.993191564438437E-8 drout = 1.631455315429714 ldrout = -1.427947792100139E-7
+ pscbe1 = 8.091529376765715E8 lpscbe1 = -2.069808714429157 pscbe2 = 1E-12
+ pvag = 0 delta = 0.01 fprout = 0
+ pdits = 0 pditsl = 0 pditsd = 0
+ lambda = 0 vtl = 0 lc = 5E-9
+ xn = 3 alpha0 = 8.506694213257144E-6 lalpha0 = -1.326670762609118E-12
+ alpha1 = 0.089171577142857 lalpha1 = 1.720506962312229E-7 beta0 = 28.332332457142854
+ lbeta0 = -2.081657060528457E-6 aigbacc = 1 bigbacc = 0
+ cigbacc = 0 nigbacc = 0 aigbinv = 0.35
+ bigbinv = 0.03 cigbinv = 6E-3 eigbinv = 1.1
+ nigbinv = 0 aigc = 0.43 bigc = 0.054
+ cigc = 0.075 aigsd = 0.43 bigsd = 0.054
+ cigsd = 0.075 dlcig = 0 nigc = 0
+ poxedge = 1 pigcd = 1 ntox = 1
+ toxref = 4.148E-9 agidl = 0 bgidl = 2.3E9
+ cgidl = 0.5 egidl = 0.8 noia = 2.5E42
+ noib = 0 noic = 0 em = 4.1E7
+ af = 1 ef = 0.84 kf = 0
+ lintnoi = -1E-7 tnoia = 1.5E7 tnoib = 9.9E6
+ ntnoi = 1 rnoia = 0.94 rnoib = 0.26
+ xpart = 0 cgso = {2.449068E-10/sw_func_tox_lv_ratio} cgdo = {2.449068E-10/sw_func_tox_lv_ratio}
+ cgbo = {1E-13/sw_func_tox_lv_ratio} ckappas = 0.6 cf = 1.4067E-12
+ clc = 1E-7 cle = 0.6 dlc = 9.87908E-9
+ dwc = 0 vfbcv = -1 noff = 3.4037
+ voffcv = -0.17287 acde = 0.4 moin = 6.9
+ cgsl = {0/sw_func_tox_lv_ratio} cgdl = {0/sw_func_tox_lv_ratio} ijthsrev = 0.1
+ ijthsfwd = 0.1 xjbvs = 1 bvs = 11.7
+ jss = 2.75E-3 jsws = 6E-10 cjs = {sw_nsd_pw_cj}
+ mjs = 0.44 mjsws = 9E-4 cjsws = {3.67354204E-11*sw_func_nsd_pw_cj}
+ cjswgs = {2.38232788E-10*sw_func_nsd_pw_cj} mjswgs = 0.8 pbs = 0.729
+ pbsws = 0.2 pbswgs = 0.95578 xrcrg1 = 12
+ xrcrg2 = 1 rbpb = 50 rbpd = 50
+ rbps = 50 rbdb = 50 rbsb = 50
+ gbmin = 1E-12 tnom = 30 ute = 1.262506997889143
+ lute = -4.819853676400192E-7 kt1 = -0.364228476514286 lkt1 = 1.640988368759452E-8
+ kt1l = 0 kt2 = -0.048405182872571 lkt2 = 1.911752584503811E-9
+ ua1 = 5.955986514324572E-9 lua1 = -1.016594662602502E-15 ub1 = -4.524249807456001E-18
+ lub1 = 8.495802448428703E-25 uc1 = -2.653294956228582E-12 luc1 = 2.096678130416571E-17
+ at = 3.525561315657149E3 lat = 5.065187629034555E-3 prt = 0
+ njs = 1.2928 xtis = 2 tpb = 1.2287E-3
+ tpbsw = 0 tpbswg = 0 tcj = 7.92E-4
+ tcjsw = 1E-5 tcjswg = 0 tvoff = 0
+ tvfbsdoff = 0 saref = 1.25E-6 sbref = 1.24E-6
+ wlod = 0 ku0 = -2.7E-8 kvsat = 0.2
+ kvth0 = 9.8E-9 tku0 = 0 llodku0 = 0
+ wlodku0 = 1 llodvth = 0 wlodvth = 1
+ lku0 = 0 wku0 = 0 pku0 = 0
+ lkvth0 = 0 wkvth0 = 2E-7 pkvth0 = 0
+ stk2 = 0 lodk2 = 1 steta0 = 0
+ lodeta0 = 1

.model nshort_model.8 nmos
+ level = 54 lmin = 1.5E-7 lmax = 1.8E-7 wmin = 7E-6
+ wmax = 1.01E-3 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 4.148E-9
+ toxm = 4.148E-9 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 9.999999999999999E22 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {2.1859E-8+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {1.1932E-8-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = 0 dwb = 0 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = 0.594819580186667 lvth0 = -1.965964275602538E-8
+ k1 = 0.819446178965333 lk1 = 1.050506912962871E-8 k2 = -0.091992990824
+ lk2 = -4.882057196623934E-9 k3 = 2 k3b = 0.54
+ w0 = 0 lpe0 = 1.0325E-7 lpeb = -7.082E-8
+ vbm = -3 dvtp0 = 0 dvtp1 = 0
+ dvt0 = 0 dvt1 = 0.53 dvt2 = -0.032
+ dvt0w = -3.58 dvt1w = 1.6706E6 dvt2w = 0.068
+ vfbsdoff = 0 u0 = 0.08215452592 lu0 = -8.197190887845112E-9
+ ua = 6.099471569173328E-9 lua = -1.072058593892447E-15 ub = -4.162341287999995E-18
+ lub = 9.026520829431672E-25 uc = 2.262880285333332E-10 luc = -2.184171335908052E-17
+ ud = 0 up = 0 lp = 1
+ eu = 1.67 vsat = 7.74854614453333E4 lvsat = 0.011033272146331
+ a0 = 1.5 ags = 1.25 b0 = 0
+ b1 = 0 keta = -0.298873933333333 lketa = 4.05375792709333E-8
+ a1 = 0 a2 = 0.42385546 rdsw = 65.968
+ rdswmin = 0 rdw = 0 rdwmin = 0
+ rsw = 0 rswmin = 0 prwb = 0
+ prwg = 0.021507 wr = 1 voff = 0.1100256
+ lvoff = -4.135817804159997E-8 voffl = 5.8197729E-9 minv = 0
+ nfactor = 10.433755181333328 lnfactor = -1.13491435899266E-6 eta0 = 0.157963749859467
+ leta0 = -1.982630242747367E-8 etab = 0.031475023122933 letab = -9.342013484634312E-9
+ dsub = 0.703398065466666 ldsub = -4.753663030570344E-8 cit = 0
+ cdsc = 0 cdscb = 0 cdscd = 0.012409066666667
+ lcdscd = -1.312958033066666E-9 pclm = 0.778108128 lpclm = -7.676865619340796E-8
+ pdiblc1 = 0.325111812096 lpdiblc1 = 7.769704881858964E-9 pdiblc2 = 5.792162294959998E-3
+ lpdiblc2 = 4.742382751629256E-10 pdiblcb = -0.449402977552439 lpdiblcb = 5.668468446307968E-8
+ drout = 1.475053670693333 ldrout = -1.183748520074542E-7 pscbe1 = 8.184366147919999E8
+ lpscbe1 = -3.519324924523709 pscbe2 = 1E-12 pvag = 0
+ delta = 0.01 fprout = 0 pdits = 0
+ pditsl = 0 pditsd = 0 lambda = 0
+ vtl = 0 lc = 5E-9 xn = 3
+ alpha0 = -7.512116426666658E-8 lalpha0 = 1.325956317594025E-14 alpha1 = 2.625266319999999
+ lalpha1 = -2.239249925395199E-7 beta0 = 19.793167999999998 lbeta0 = -7.483860788479997E-7
+ aigbacc = 1 bigbacc = 0 cigbacc = 0
+ nigbacc = 0 aigbinv = 0.35 bigbinv = 0.03
+ cigbinv = 6E-3 eigbinv = 1.1 nigbinv = 0
+ aigc = 0.43 bigc = 0.054 cigc = 0.075
+ aigsd = 0.43 bigsd = 0.054 cigsd = 0.075
+ dlcig = 0 nigc = 0 poxedge = 1
+ pigcd = 1 ntox = 1 toxref = 4.148E-9
+ agidl = 0 bgidl = 2.3E9 cgidl = 0.5
+ egidl = 0.8 noia = 2.5E42 noib = 0
+ noic = 0 em = 4.1E7 af = 1
+ ef = 0.84 kf = 0 lintnoi = -1E-7
+ tnoia = 1.5E7 tnoib = 9.9E6 ntnoi = 1
+ rnoia = 0.94 rnoib = 0.26 xpart = 0
+ cgso = {2.449068E-10/sw_func_tox_lv_ratio} cgdo = {2.449068E-10/sw_func_tox_lv_ratio} cgbo = {1E-13/sw_func_tox_lv_ratio}
+ ckappas = 0.6 cf = 1.4067E-12 clc = 1E-7
+ cle = 0.6 dlc = 9.87908E-9 dwc = 0
+ vfbcv = -1 noff = 3.4037 voffcv = -0.17287
+ acde = 0.4 moin = 6.9 cgsl = {0/sw_func_tox_lv_ratio}
+ cgdl = {0/sw_func_tox_lv_ratio} ijthsrev = 0.1 ijthsfwd = 0.1
+ xjbvs = 1 bvs = 11.7 jss = 2.75E-3
+ jsws = 6E-10 cjs = {sw_nsd_pw_cj} mjs = 0.44
+ mjsws = 9E-4 cjsws = {3.67354204E-11*sw_func_nsd_pw_cj} cjswgs = {2.38232788E-10*sw_func_nsd_pw_cj}
+ mjswgs = 0.8 pbs = 0.729 pbsws = 0.2
+ pbswgs = 0.95578 xrcrg1 = 12 xrcrg2 = 1
+ rbpb = 50 rbpd = 50 rbps = 50
+ rbdb = 50 rbsb = 50 gbmin = 1E-12
+ tnom = 30 ute = -9.495419167253328 lute = 1.197714192080666E-6
+ kt1 = -0.442902553381333 lkt1 = 2.869373935330785E-8 kt1l = 0
+ kt2 = -0.0644473841808 lkt2 = 4.416517727965387E-9 ua1 = -1.123856160673066E-8
+ lua1 = 1.668093302826578E-15 ub1 = 7.039606710197328E-18 lub1 = -9.559540563974501E-25
+ uc1 = 1.73590446640001E-11 luc1 = 1.784213464522168E-17 at = 4.957831755386664E4
+ lat = -2.125305518974522E-3 prt = 0 njs = 1.2928
+ xtis = 2 tpb = 1.2287E-3 tpbsw = 0
+ tpbswg = 0 tcj = 7.92E-4 tcjsw = 1E-5
+ tcjswg = 0 tvoff = 0 tvfbsdoff = 0
+ saref = 1.1E-6 sbref = 1.1E-6 wlod = 0
+ ku0 = -2.7E-8 kvsat = 0.2 kvth0 = 9.8E-9
+ tku0 = 0 llodku0 = 0 wlodku0 = 1
+ llodvth = 0 wlodvth = 1 lku0 = 0
+ wku0 = 0 pku0 = 0 lkvth0 = 0
+ wkvth0 = 2E-7 pkvth0 = 0 stk2 = 0
+ lodk2 = 1 steta0 = 0 lodeta0 = 1

.model nshort_model.9 nmos
+ level = 54 lmin = 8E-6 lmax = 2.02E-5 wmin = 5E-6
+ wmax = 7E-6 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 4.148E-9
+ toxm = 4.148E-9 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 9.999999999999999E22 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {2.1859E-8+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {1.1932E-8-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = 0 dwb = 0 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = 0.5187147 k1 = 0.53705506214712
+ wk1 = 2.650752369040756E-8 k2 = -0.02665245231549 wk2 = -5.018170325606322E-10
+ k3 = 2 k3b = 0.54 w0 = 0
+ lpe0 = 1.0325E-7 lpeb = -7.082E-8 vbm = -3
+ dvtp0 = 0 dvtp1 = 0 dvt0 = 0
+ dvt1 = 0.53 dvt2 = -0.032 dvt0w = -3.58
+ dvt1w = 1.6706E6 dvt2w = 0.068 vfbsdoff = 0
+ u0 = 0.0330727153208 wu0 = -8.426250962405228E-9 ua = -8.483379519471496E-10
+ wua = 6.238002890000825E-16 ub = 1.886474514342E-18 wub = -1.476697033431996E-24
+ uc = 5.533574871900001E-11 wuc = -4.23898345265028E-17 ud = 0
+ up = 0 lp = 1 eu = 1.67
+ vsat = 8E4 a0 = 1.2750373037511 wa0 = 4.144670811456904E-7
+ ags = 0.4171236043699 wags = -8.315751231085662E-8 b0 = 0
+ b1 = 7.329634002478404E-24 wb1 = -3.632773307307167E-29 keta = -0.015256722396137
+ wketa = 4.495234570604608E-8 a1 = 0 a2 = 0.42385546
+ rdsw = 65.968 rdswmin = 0 rdw = 0
+ rdwmin = 0 rsw = 0 rswmin = 0
+ prwb = 0 prwg = 0.021507 wr = 1
+ voff = -0.10821273063364 wvoff = 2.048020293243856E-8 voffl = 5.8197729E-9
+ minv = 0 nfactor = 2.43689254434 wnfactor = 1.366335211293459E-6
+ eta0 = 0.08 etab = -0.07 dsub = 0.56
+ cit = 0 cdsc = 0 cdscb = 0
+ cdscd = 5.4E-3 pclm = -0.098993677806 wpclm = 8.716894561476778E-7
+ pdiblc1 = 0.39 pdiblc2 = 2.7755113119418E-3 wpdiblc2 = 2.07260605249627E-9
+ pdiblcb = -0.025 drout = 0.56 pscbe1 = 9.037191253642601E8
+ wpscbe1 = -1.036798809754026E3 pscbe2 = 1E-12 pvag = 0
+ delta = 0.01 fprout = 0 pdits = 0
+ pditsl = 0 pditsd = 0 lambda = 0
+ vtl = 0 lc = 5E-9 xn = 3
+ alpha0 = 3E-8 alpha1 = 0.85 beta0 = 13.86
+ aigbacc = 1 bigbacc = 0 cigbacc = 0
+ nigbacc = 0 aigbinv = 0.35 bigbinv = 0.03
+ cigbinv = 6E-3 eigbinv = 1.1 nigbinv = 0
+ aigc = 0.43 bigc = 0.054 cigc = 0.075
+ aigsd = 0.43 bigsd = 0.054 cigsd = 0.075
+ dlcig = 0 nigc = 0 poxedge = 1
+ pigcd = 1 ntox = 1 toxref = 4.148E-9
+ agidl = 0 bgidl = 2.3E9 cgidl = 0.5
+ egidl = 0.8 noia = 2.5E42 noib = 0
+ noic = 0 em = 4.1E7 af = 1
+ ef = 0.84 kf = 0 lintnoi = -1E-7
+ tnoia = 1.5E7 tnoib = 9.9E6 ntnoi = 1
+ rnoia = 0.94 rnoib = 0.26 xpart = 0
+ cgso = {2.449068E-10/sw_func_tox_lv_ratio} cgdo = {2.449068E-10/sw_func_tox_lv_ratio} cgbo = {1E-13/sw_func_tox_lv_ratio}
+ ckappas = 0.6 cf = 1.4067E-12 clc = 1E-7
+ cle = 0.6 dlc = 9.87908E-9 dwc = 0
+ vfbcv = -1 noff = 3.4037 voffcv = -0.17287
+ acde = 0.4 moin = 6.9 cgsl = {0/sw_func_tox_lv_ratio}
+ cgdl = {0/sw_func_tox_lv_ratio} ijthsrev = 0.1 ijthsfwd = 0.1
+ xjbvs = 1 bvs = 11.7 jss = 2.75E-3
+ jsws = 6E-10 cjs = {sw_nsd_pw_cj} mjs = 0.44
+ mjsws = 9E-4 cjsws = {3.67354204E-11*sw_func_nsd_pw_cj} cjswgs = {2.38232788E-10*sw_func_nsd_pw_cj}
+ mjswgs = 0.8 pbs = 0.729 pbsws = 0.2
+ pbswgs = 0.95578 xrcrg1 = 12 xrcrg2 = 1
+ rbpb = 50 rbpd = 50 rbps = 50
+ rbdb = 50 rbsb = 50 gbmin = 1E-12
+ tnom = 30 ute = -1.6391866877 wute = -1.21187692851287E-6
+ kt1 = -0.28485353683 wkt1 = -1.960034235731348E-7 kt1l = 0
+ kt2 = -0.044827209992594 wkt2 = -3.381636551332185E-9 ua1 = 6.657642457200001E-10
+ wua1 = -2.015542681105614E-15 ub1 = -9.909460495700003E-19 wub1 = 2.4439230747549E-24
+ uc1 = 1.2862847900826E-11 wuc1 = 2.063835028581233E-17 at = 1.4E5
+ prt = 0 njs = 1.2928 xtis = 2
+ tpb = 1.2287E-3 tpbsw = 0 tpbswg = 0
+ tcj = 7.92E-4 tcjsw = 1E-5 tcjswg = 0
+ tvoff = 0 tvfbsdoff = 0 saref = 3E-6
+ sbref = 3E-6 wlod = 0 ku0 = -2.7E-8
+ kvsat = 0.2 kvth0 = 9.8E-9 tku0 = 0
+ llodku0 = 0 wlodku0 = 1 llodvth = 0
+ wlodvth = 1 lku0 = 0 wku0 = 0
+ pku0 = 0 lkvth0 = 0 wkvth0 = 2E-7
+ pkvth0 = 0 stk2 = 0 lodk2 = 1
+ steta0 = 0 lodeta0 = 1

.model nshort_model.10 nmos
+ level = 54 lmin = 4E-6 lmax = 8E-6 wmin = 5E-6
+ wmax = 7E-6 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 4.148E-9
+ toxm = 4.148E-9 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 9.999999999999999E22 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {2.1859E-8+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {1.1932E-8-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = 0 dwb = 0 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = 0.514861965187682 lvth0 = 3.890276704946321E-8
+ wvth0 = -1.422559662518131E-8 pvth0 = 7.295844208250089E-14 k1 = 0.524711243807652
+ lk1 = 9.845597383489342E-8 wk1 = 4.912095597296223E-8 pk1 = -1.803678113124465E-13
+ k2 = -0.019213029200116 lk2 = -5.933785052977059E-8 wk2 = -1.115997734504156E-8
+ pk2 = 8.501093616215041E-14 k3 = 2 k3b = 0.54
+ w0 = 0 lpe0 = 1.0325E-7 lpeb = -7.082E-8
+ vbm = -3 dvtp0 = 0 dvtp1 = 0
+ dvt0 = 0 dvt1 = 0.53 dvt2 = -0.032
+ dvt0w = -3.58 dvt1w = 1.6706E6 dvt2w = 0.068
+ vfbsdoff = 0 u0 = 0.034470037136056 lu0 = -1.114522883425205E-8
+ wu0 = -1.59454408185693E-8 pu0 = 5.997408090258504E-14 ua = -8.875308152487672E-10
+ lua = 3.126076079231105E-16 wua = 8.606698489748808E-16 pua = -1.889303824619149E-21
+ ub = 2.069398669602868E-18 lub = -1.459027940045796E-24 wub = -2.553784995143585E-24
+ pub = 8.591000066574424E-30 uc = 1.754519486956829E-10 luc = -9.580631468172194E-16
+ wuc = -8.340638804580831E-16 puc = 6.314499858020532E-21 ud = 0
+ up = 0 lp = 1 eu = 1.67
+ vsat = 8E4 a0 = 1.649897199300823 la0 = -2.989933507850385E-6
+ wa0 = -1.530071155902545E-6 pa0 = 1.550990143589697E-11 ags = 0.531557742938164
+ lags = -9.127422522633187E-7 wags = -9.678943845638612E-7 pags = 7.056781617304592E-12
+ b0 = 0 b1 = 1.461553940849802E-23 lb1 = -5.811337240154769E-29
+ wb1 = -7.24387348906294E-29 pb1 = 2.880262615930876E-34 keta = -0.028499150973664
+ lketa = 1.056234113046414E-7 wketa = 8.996208595294972E-8 pketa = -3.59003809533977E-13
+ a1 = 0 a2 = 0.42385546 rdsw = 65.968
+ rdswmin = 0 rdw = 0 rdwmin = 0
+ rsw = 0 rswmin = 0 prwb = 0
+ prwg = 0.021507 wr = 1 voff = -0.117643830538068
+ lvoff = 7.522373546730369E-8 wvoff = 6.10572676628412E-8 pvoff = -3.236481867704948E-13
+ voffl = 5.8197729E-9 minv = 0 nfactor = 2.199884559689013
+ lnfactor = 1.890407918662182E-6 wnfactor = 2.730002323311536E-6 pnfactor = -1.087679434418342E-11
+ eta0 = 0.08 etab = -0.07 dsub = 0.56
+ cit = 0 cdsc = 0 cdscb = 0
+ cdscd = 5.4E-3 pclm = -1.019244330754529 lpclm = 7.34004436200627E-6
+ wpclm = 3.396067242954099E-6 ppclm = -2.013478054294703E-11 pdiblc1 = 0.39
+ pdiblc2 = 2.814622144645338E-3 lpdiblc2 = -3.11953320716663E-10 wpdiblc2 = 1.682108545390056E-9
+ ppdiblc2 = 3.114661224340133E-15 pdiblcb = -0.025 drout = 0.56
+ pscbe1 = 1.004186824163253E9 lpscbe1 = -801.344029227806 wpscbe1 = -2.04909870364525E3
+ ppscbe1 = 8.07424162646197E-3 pscbe2 = 1E-12 pvag = 0
+ delta = 0.01 fprout = 0 pdits = 0
+ pditsl = 0 pditsd = 0 lambda = 0
+ vtl = 0 lc = 5E-9 xn = 3
+ alpha0 = 3E-8 alpha1 = 0.85 beta0 = 13.86
+ aigbacc = 1 bigbacc = 0 cigbacc = 0
+ nigbacc = 0 aigbinv = 0.35 bigbinv = 0.03
+ cigbinv = 6E-3 eigbinv = 1.1 nigbinv = 0
+ aigc = 0.43 bigc = 0.054 cigc = 0.075
+ aigsd = 0.43 bigsd = 0.054 cigsd = 0.075
+ dlcig = 0 nigc = 0 poxedge = 1
+ pigcd = 1 ntox = 1 toxref = 4.148E-9
+ agidl = 0 bgidl = 2.3E9 cgidl = 0.5
+ egidl = 0.8 noia = 2.5E42 noib = 0
+ noic = 0 em = 4.1E7 af = 1
+ ef = 0.84 kf = 0 lintnoi = -1E-7
+ tnoia = 1.5E7 tnoib = 9.9E6 ntnoi = 1
+ rnoia = 0.94 rnoib = 0.26 xpart = 0
+ cgso = {2.449068E-10/sw_func_tox_lv_ratio} cgdo = {2.449068E-10/sw_func_tox_lv_ratio} cgbo = {1E-13/sw_func_tox_lv_ratio}
+ ckappas = 0.6 cf = 1.4067E-12 clc = 1E-7
+ cle = 0.6 dlc = 9.87908E-9 dwc = 0
+ vfbcv = -1 noff = 3.4037 voffcv = -0.17287
+ acde = 0.4 moin = 6.9 cgsl = {0/sw_func_tox_lv_ratio}
+ cgdl = {0/sw_func_tox_lv_ratio} ijthsrev = 0.1 ijthsfwd = 0.1
+ xjbvs = 1 bvs = 11.7 jss = 2.75E-3
+ jsws = 6E-10 cjs = {sw_nsd_pw_cj} mjs = 0.44
+ mjsws = 9E-4 cjsws = {3.67354204E-11*sw_func_nsd_pw_cj} cjswgs = {2.38232788E-10*sw_func_nsd_pw_cj}
+ mjswgs = 0.8 pbs = 0.729 pbsws = 0.2
+ pbswgs = 0.95578 xrcrg1 = 12 xrcrg2 = 1
+ rbpb = 50 rbpd = 50 rbps = 50
+ rbdb = 50 rbsb = 50 gbmin = 1E-12
+ tnom = 30 ute = -1.119515970036249 lute = -4.144964319303681E-6
+ wute = -4.5516447110251E-6 pute = 2.663844204173598E-11 kt1 = -0.25967447552086
+ lkt1 = -2.00831617354038E-7 wkt1 = -3.565658870012505E-7 pkt1 = 1.280668044797677E-12
+ kt1l = 0 kt2 = -0.03215028598288 lkt2 = -1.011128699631404E-7
+ wkt2 = -8.381152134652494E-8 pkt2 = 6.415196995907897E-13 ua1 = 1.9194868601037E-9
+ lua1 = -9.999862078599947E-15 wua1 = -9.374855505915913E-15 pua1 = 5.869887995723112E-20
+ ub1 = -2.193186578214897E-18 lub1 = 9.589233961183593E-24 wub1 = 9.024070988991411E-24
+ pub1 = -5.248415466406676E-29 uc1 = -2.774183418740579E-11 luc1 = 3.238684665725007E-16
+ wuc1 = 2.026400665814326E-16 puc1 = -1.451670441407283E-21 at = 1.4E5
+ prt = 0 njs = 1.2928 xtis = 2
+ tpb = 1.2287E-3 tpbsw = 0 tpbswg = 0
+ tcj = 7.92E-4 tcjsw = 1E-5 tcjswg = 0
+ tvoff = 0 tvfbsdoff = 0 saref = 3E-6
+ sbref = 3E-6 wlod = 0 ku0 = -2.7E-8
+ kvsat = 0.2 kvth0 = 9.8E-9 tku0 = 0
+ llodku0 = 0 wlodku0 = 1 llodvth = 0
+ wlodvth = 1 lku0 = 0 wku0 = 0
+ pku0 = 0 lkvth0 = 0 wkvth0 = 2E-7
+ pkvth0 = 0 stk2 = 0 lodk2 = 1
+ steta0 = 0 lodeta0 = 1

.model nshort_model.11 nmos
+ level = 54 lmin = 2E-6 lmax = 4E-6 wmin = 5E-6
+ wmax = 7E-6 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 4.148E-9
+ toxm = 4.148E-9 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 9.999999999999999E22 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {2.1859E-8+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {1.1932E-8-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = 0 dwb = 0 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = 0.51690684343716 lvth0 = 3.077205302609519E-8
+ wvth0 = 1.14135897192752E-8 pvth0 = -2.898644975240104E-14 k1 = 0.575533903540702
+ lk1 = -1.036218331454398E-7 wk1 = -1.766487393951152E-7 pk1 = 7.173232021495994E-13
+ k2 = -0.043352844857489 lk2 = 3.664533953887408E-8 wk2 = 8.385648890813032E-8
+ pk2 = -2.927874558998715E-13 k3 = 2 k3b = 0.54
+ w0 = 0 lpe0 = 1.0325E-7 lpeb = -7.082E-8
+ vbm = -3 dvtp0 = 0 dvtp1 = 0
+ dvt0 = 0 dvt1 = 0.53 dvt2 = -0.032
+ dvt0w = -3.58 dvt1w = 1.6706E6 dvt2w = 0.068
+ vfbsdoff = 0 u0 = 0.033383605099746 lu0 = -6.82542730312602E-9
+ wu0 = -1.229844233093496E-9 pu0 = 1.462867557597635E-15 ua = -4.089115672306983E-10
+ lua = -1.590447614414462E-15 wua = -1.212818207960921E-15 pua = 6.355166684133342E-21
+ ub = 1.219303834670351E-18 lub = 1.921064736543442E-24 wub = 2.118126315932818E-24
+ pub = -9.985154686203658E-30 uc = -2.097160149949759E-10 luc = 5.734170596599017E-16
+ wuc = 1.541281883502334E-15 puc = -3.130197946509985E-21 ud = 0
+ up = 0 lp = 1 eu = 1.67
+ vsat = 8E4 a0 = 0.506713346936195 la0 = 1.555520962155299E-6
+ wa0 = 5.169582504252088E-6 pa0 = -1.112883266977564E-11 ags = 0.01121682116155
+ lags = 1.156204019085862E-6 wags = 1.690610240424994E-6 pags = -3.513794328280096E-12
+ b0 = 0 b1 = 0 keta = -1.528191735747104E-5
+ lketa = -7.63232586942559E-9 wketa = -2.642739692980208E-8 pketa = 1.037766033775162E-13
+ a1 = 0 a2 = 0.42385546 rdsw = 65.968
+ rdswmin = 0 rdw = 0 rdwmin = 0
+ rsw = 0 rswmin = 0 prwb = 0
+ prwg = 0.021507 wr = 1 voff = -0.088721265394765
+ lvoff = -3.977631701132865E-8 wvoff = -8.808335946553013E-8 pvoff = 2.693552298171991E-13
+ voffl = 5.8197729E-9 minv = 0 nfactor = 2.672677675829692
+ lnfactor = 1.051818902304774E-8 wnfactor = -5.449500865560848E-7 pnfactor = 2.144861830977985E-12
+ eta0 = 0.158551406 leta0 = -3.123310732472159E-7 etab = -0.138668351310661
+ letab = 2.73034703706968E-7 wetab = -1.176909133861078E-11 petab = 4.679550775873851E-17
+ dsub = 0.8564204 ldsub = -1.1786078235744E-6 cit = 0
+ cdsc = 0 cdscb = 0 cdscd = 5.4E-3
+ pclm = 0.834777993773728 lpclm = -3.180054735421614E-8 wpclm = -1.531916168788979E-6
+ ppclm = -5.404482921125471E-13 pdiblc1 = 0.39 pdiblc2 = 1.32990405975453E-3
+ lpdiblc2 = 5.591487706468735E-9 wpdiblc2 = 4.126490088005316E-10 ppdiblc2 = 8.162204988317059E-15
+ pdiblcb = -0.025 drout = 0.56 pscbe1 = 8.052652765266876E8
+ lpscbe1 = -10.404902494342187 wpscbe1 = -36.62674832761898 ppscbe1 = 7.237943593314765E-5
+ pscbe2 = 1E-12 pvag = 0 delta = 0.01
+ fprout = 0 pdits = 0 pditsl = 0
+ pditsd = 0 lambda = 0 vtl = 0
+ lc = 5E-9 xn = 3 alpha0 = 3E-8
+ alpha1 = 0.85 beta0 = 13.86 aigbacc = 1
+ bigbacc = 0 cigbacc = 0 nigbacc = 0
+ aigbinv = 0.35 bigbinv = 0.03 cigbinv = 6E-3
+ eigbinv = 1.1 nigbinv = 0 aigc = 0.43
+ bigc = 0.054 cigc = 0.075 aigsd = 0.43
+ bigsd = 0.054 cigsd = 0.075 dlcig = 0
+ nigc = 0 poxedge = 1 pigcd = 1
+ ntox = 1 toxref = 4.148E-9 agidl = 0
+ bgidl = 2.3E9 cgidl = 0.5 egidl = 0.8
+ noia = 2.5E42 noib = 0 noic = 0
+ em = 4.1E7 af = 1 ef = 0.84
+ kf = 0 lintnoi = -1E-7 tnoia = 1.5E7
+ tnoib = 9.9E6 ntnoi = 1 rnoia = 0.94
+ rnoib = 0.26 xpart = 0 cgso = {2.449068E-10/sw_func_tox_lv_ratio}
+ cgdo = {2.449068E-10/sw_func_tox_lv_ratio} cgbo = {1E-13/sw_func_tox_lv_ratio} ckappas = 0.6
+ cf = 1.4067E-12 clc = 1E-7 cle = 0.6
+ dlc = 9.87908E-9 dwc = 0 vfbcv = -1
+ noff = 3.4037 voffcv = -0.17287 acde = 0.4
+ moin = 6.9 cgsl = {0/sw_func_tox_lv_ratio} cgdl = {0/sw_func_tox_lv_ratio}
+ ijthsrev = 0.1 ijthsfwd = 0.1 xjbvs = 1
+ bvs = 11.7 jss = 2.75E-3 jsws = 6E-10
+ cjs = {sw_nsd_pw_cj} mjs = 0.44 mjsws = 9E-4
+ cjsws = {3.67354204E-11*sw_func_nsd_pw_cj} cjswgs = {2.38232788E-10*sw_func_nsd_pw_cj} mjswgs = 0.8
+ pbs = 0.729 pbsws = 0.2 pbswgs = 0.95578
+ xrcrg1 = 12 xrcrg2 = 1 rbpb = 50
+ rbpd = 50 rbps = 50 rbdb = 50
+ rbsb = 50 gbmin = 1E-12 tnom = 30
+ ute = -2.533689067872448 lute = 1.477980245234353E-6 wute = 3.783099279386647E-6
+ pute = -6.501633589323831E-12 kt1 = -0.304681311684496 lkt1 = -2.187831583770234E-8
+ wkt1 = -1.199379322707409E-8 pkt1 = -8.939746185320198E-14 kt1l = 0
+ kt2 = -0.058147650511164 lkt2 = 2.256187042891775E-9 wkt2 = 8.157323401053458E-8
+ pkt2 = -1.607258003560759E-14 ua1 = -1.721514168753613E-9 lua1 = 4.477253188276655E-15
+ wua1 = 1.111578179065378E-14 pua1 = -2.27746806606023E-20 ub1 = 1.23986714426398E-18
+ lub1 = -4.061054534698681E-24 wub1 = -1.00190435314664E-23 pub1 = 2.32338585328483E-29
+ uc1 = 6.727091943573324E-11 luc1 = -5.391516356759274E-17 wuc1 = -2.985607599961264E-16
+ puc1 = 5.411722083775055E-22 at = 1.677727274205532E5 lat = -0.110428141315049
+ wat = -0.02095053598851 pat = 8.33021803632117E-8 prt = 0
+ njs = 1.2928 xtis = 2 tpb = 1.2287E-3
+ tpbsw = 0 tpbswg = 0 tcj = 7.92E-4
+ tcjsw = 1E-5 tcjswg = 0 tvoff = 0
+ tvfbsdoff = 0 saref = 3E-6 sbref = 3E-6
+ wlod = 0 ku0 = -2.7E-8 kvsat = 0.2
+ kvth0 = 9.8E-9 tku0 = 0 llodku0 = 0
+ wlodku0 = 1 llodvth = 0 wlodvth = 1
+ lku0 = 0 wku0 = 0 pku0 = 0
+ lkvth0 = 0 wkvth0 = 2E-7 pkvth0 = 0
+ stk2 = 0 lodk2 = 1 steta0 = 0
+ lodeta0 = 1

.model nshort_model.12 nmos
+ level = 54 lmin = 1E-6 lmax = 2E-6 wmin = 5E-6
+ wmax = 7E-6 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 4.148E-9
+ toxm = 4.148E-9 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 9.999999999999999E22 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {2.1859E-8+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {1.1932E-8-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = 0 dwb = 0 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = 0.514368709462509 lvth0 = 3.578775094622736E-8
+ wvth0 = -4.367374610919243E-8 pvth0 = 7.987361772232366E-14 k1 = 0.434089457827375
+ lk1 = 1.758916280287128E-7 wk1 = 5.763314290519126E-7 pk1 = -7.706680160046362E-13
+ k2 = 0.010291856684145 lk2 = -6.936388638680422E-8 wk2 = -2.186303862509402E-7
+ pk2 = 3.049677476294735E-13 k3 = 2 k3b = 0.54
+ w0 = 0 lpe0 = 1.0325E-7 lpeb = -7.082E-8
+ vbm = -3 dvtp0 = 0 dvtp1 = 0
+ dvt0 = 0 dvt1 = 0.53 dvt2 = -0.032
+ dvt0w = -3.58 dvt1w = 1.6706E6 dvt2w = 0.068
+ vfbsdoff = 0 u0 = 0.03384188646021 lu0 = -7.731053597666928E-9
+ wu0 = -8.932636691687881E-10 pu0 = 7.977385883257185E-16 ua = -9.299748179488245E-10
+ lua = -5.60755766393347E-16 wua = 3.545575809160351E-15 pua = -3.048067035284618E-21
+ ub = 2.074615849962149E-18 lub = 2.308518718927696E-25 wub = -5.362545924103436E-24
+ pub = 4.797671031532622E-30 uc = 7.461009665150011E-11 luc = 1.154999469528129E-17
+ wuc = 8.920838519876666E-17 puc = -2.607032318663673E-22 ud = 0
+ up = 0 lp = 1 eu = 1.67
+ vsat = 2.043538776733193E4 lvsat = 0.117707774559016 wvsat = 0.276505610998143
+ pvsat = -5.464126920954264E-7 a0 = 2.240715044656126 la0 = -1.871102216770174E-6
+ wa0 = -6.089017015773056E-6 pa0 = 1.111969115132877E-11 ags = 1.178946724951263
+ lags = -1.151389082069527E-6 wags = -6.244912459396909E-6 pags = 1.216787775765516E-11
+ b0 = 0 b1 = 0 keta = 0.051445067799949
+ lketa = -1.093249755183855E-7 wketa = 8.223904274173894E-8 pketa = -1.109630600492442E-13
+ a1 = 0 a2 = 0.42385546 rdsw = 65.968
+ rdswmin = 0 rdw = 0 rdwmin = 0
+ rsw = 0 rswmin = 0 prwb = 0
+ prwg = 0.021507 wr = 1 voff = -0.10407400415042
+ lvoff = -9.43721725768379E-9 wvoff = 1.42104150412363E-7 pvoff = -1.85526595202861E-13
+ voffl = 5.8197729E-9 minv = 0 nfactor = 2.605050779692767
+ lnfactor = 1.441581330474852E-7 wnfactor = 1.834306897719281E-6 pnfactor = -2.556873548899999E-12
+ eta0 = -6.411041806166857E-3 leta0 = 1.365715851067135E-8 weta0 = 3.428240497958349E-8
+ peta0 = -6.77466946467342E-14 etab = -9.63205325672294E-4 letab = 9.10607340775536E-10
+ wetab = 1.939510043361299E-9 petab = -3.809197436370392E-15 dsub = 1.133108040820545
+ ldsub = -1.725380231354949E-6 wdsub = -6.073585748415222E-6 pdsub = 1.200223144653026E-11
+ cit = 0 cdsc = 0 cdscb = 0
+ cdscd = 5.4E-3 pclm = 1.096795738110111 lpclm = -5.495832445761399E-7
+ wpclm = -2.602847633246711E-6 ppclm = 1.575857928335097E-12 pdiblc1 = -0.188441663672555
+ lpdiblc1 = 1.143079395483228E-6 wpdiblc1 = 1.870182013222829E-6 ppdiblc1 = -3.695734002882108E-12
+ pdiblc2 = 6.815002986727553E-3 lpdiblc2 = -5.247813746684025E-9 wpdiblc2 = -8.490490509427675E-9
+ ppdiblc2 = 2.575601950331047E-14 pdiblcb = -0.048987242130015 lpdiblcb = 4.740205271384014E-8
+ wpdiblcb = -1.593947539938265E-9 ppdiblcb = 3.149857115783443E-15 drout = 0.8528408
+ ldrout = -5.786932471488001E-7 pscbe1 = 2.326916344252413E9 lpscbe1 = -3.017394356865586E3
+ wpscbe1 = -6.962207506759606E3 ppscbe1 = 0.013758268893578 pscbe2 = 1E-12
+ pvag = 0 delta = 0.01 fprout = 0
+ pdits = 0 pditsl = 0 pditsd = 0
+ lambda = 0 vtl = 0 lc = 5E-9
+ xn = 3 alpha0 = 3.850882118112005E-7 lalpha0 = -7.017025985357398E-13
+ walpha0 = -2.019271745361316E-11 palpha0 = 3.99035558979133E-17 alpha1 = 0.816811376
+ lalpha1 = 6.558523467686407E-8 beta0 = 11.824214740159743 lbeta0 = 4.022988540239684E-6
+ wbeta0 = -4.661152278875665E-6 pbeta0 = 9.21107081976824E-12 aigbacc = 1
+ bigbacc = 0 cigbacc = 0 nigbacc = 0
+ aigbinv = 0.35 bigbinv = 0.03 cigbinv = 6E-3
+ eigbinv = 1.1 nigbinv = 0 aigc = 0.43
+ bigc = 0.054 cigc = 0.075 aigsd = 0.43
+ bigsd = 0.054 cigsd = 0.075 dlcig = 0
+ nigc = 0 poxedge = 1 pigcd = 1
+ ntox = 1 toxref = 4.148E-9 agidl = 0
+ bgidl = 2.3E9 cgidl = 0.5 egidl = 0.8
+ noia = 2.5E42 noib = 0 noic = 0
+ em = 4.1E7 af = 1 ef = 0.84
+ kf = 0 lintnoi = -1E-7 tnoia = 1.5E7
+ tnoib = 9.9E6 ntnoi = 1 rnoia = 0.94
+ rnoib = 0.26 xpart = 0 cgso = {2.449068E-10/sw_func_tox_lv_ratio}
+ cgdo = {2.449068E-10/sw_func_tox_lv_ratio} cgbo = {1E-13/sw_func_tox_lv_ratio} ckappas = 0.6
+ cf = 1.4067E-12 clc = 1E-7 cle = 0.6
+ dlc = 9.87908E-9 dwc = 0 vfbcv = -1
+ noff = 3.4037 voffcv = -0.17287 acde = 0.4
+ moin = 6.9 cgsl = {0/sw_func_tox_lv_ratio} cgdl = {0/sw_func_tox_lv_ratio}
+ ijthsrev = 0.1 ijthsfwd = 0.1 xjbvs = 1
+ bvs = 11.7 jss = 2.75E-3 jsws = 6E-10
+ cjs = {sw_nsd_pw_cj} mjs = 0.44 mjsws = 9E-4
+ cjsws = {3.67354204E-11*sw_func_nsd_pw_cj} cjswgs = {2.38232788E-10*sw_func_nsd_pw_cj} mjswgs = 0.8
+ pbs = 0.729 pbsws = 0.2 pbswgs = 0.95578
+ xrcrg1 = 12 xrcrg2 = 1 rbpb = 50
+ rbpd = 50 rbps = 50 rbdb = 50
+ rbsb = 50 gbmin = 1E-12 tnom = 30
+ ute = -2.561971268216158 lute = 1.533869719492769E-6 wute = 2.695685041105775E-7
+ pute = 4.415810628071198E-13 kt1 = -0.359948466175884 lkt1 = 8.73370977702914E-8
+ wkt1 = -9.806652819008198E-8 pkt1 = 8.069396832565656E-14 kt1l = 0
+ kt2 = -0.08698809059532 lkt2 = 5.924881894903557E-8 wkt2 = 1.457790957302304E-7
+ pkt2 = -1.429520947909204E-13 ua1 = -8.561527014636378E-10 lua1 = 2.767181239752113E-15
+ wua1 = -2.339774546732115E-15 pua1 = 3.815328617734101E-21 ub1 = -3.464362798299158E-19
+ lub1 = -9.263032314234665E-25 wub1 = 4.605306502872922E-24 pub1 = -5.665846046610872E-30
+ uc1 = 1.17750393204133E-11 luc1 = 5.575224297997512E-17 wuc1 = 3.960554356093764E-17
+ puc1 = -1.270903980685366E-22 at = 1.562147447217006E5 lat = -0.087587995616469
+ wat = 0.063082997004157 pat = -8.27595093907865E-8 prt = 0
+ njs = 1.2928 xtis = 2 tpb = 1.2287E-3
+ tpbsw = 0 tpbswg = 0 tcj = 7.92E-4
+ tcjsw = 1E-5 tcjswg = 0 tvoff = 0
+ tvfbsdoff = 0 saref = 3E-6 sbref = 3E-6
+ wlod = 0 ku0 = -2.7E-8 kvsat = 0.2
+ kvth0 = 9.8E-9 tku0 = 0 llodku0 = 0
+ wlodku0 = 1 llodvth = 0 wlodvth = 1
+ lku0 = 0 wku0 = 0 pku0 = 0
+ lkvth0 = 0 wkvth0 = 2E-7 pkvth0 = 0
+ stk2 = 0 lodk2 = 1 steta0 = 0
+ lodeta0 = 1

.model nshort_model.13 nmos
+ level = 54 lmin = 5E-7 lmax = 1E-6 wmin = 5E-6
+ wmax = 7E-6 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 4.148E-9
+ toxm = 4.148E-9 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 9.999999999999999E22 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {2.1859E-8+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {1.1932E-8-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = 0 dwb = 0 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = 0.541070442633641 lvth0 = 9.723227935491056E-9
+ wvth0 = -1.990202567734794E-8 pvth0 = 5.66691856268647E-14 k1 = 0.71742673412354
+ lk1 = -1.006840875059212E-7 wk1 = -2.822257427043878E-7 pk1 = 6.740054740487191E-14
+ k2 = -0.106360861512381 lk2 = 4.450503134268032E-8 wk2 = 1.547920099728853E-7
+ pk2 = -5.954329653086669E-14 k3 = 2 k3b = 0.54
+ w0 = 0 lpe0 = 1.0325E-7 lpeb = -7.082E-8
+ vbm = -3 dvtp0 = 0 dvtp1 = 0
+ dvt0 = 0 dvt1 = 0.53 dvt2 = -0.032
+ dvt0w = -3.58 dvt1w = 1.6706E6 dvt2w = 0.068
+ vfbsdoff = 0 u0 = 0.029104774260518 lu0 = -3.106987843508501E-9
+ wu0 = -7.266506832111083E-9 pu0 = 7.018890676427559E-15 ua = -1.278540519869651E-9
+ lua = -2.20508236383159E-16 wua = -6.451937388303618E-17 pua = 4.758768363106218E-22
+ ub = 2.255126143608551E-18 lub = 5.464927589394545E-26 wub = -1.969794007794512E-25
+ pub = -2.44624412278759E-31 uc = 8.709476102894867E-11 luc = -6.36735651463838E-19
+ wuc = -3.273185510544497E-16 puc = 1.458837055801024E-22 ud = 0
+ up = 0 lp = 1 eu = 1.67
+ vsat = 1.852060169569901E5 lvsat = -0.04313076833566 wvsat = -0.679433208277503
+ pvsat = 3.867136031970258E-7 a0 = -0.796127191879444 la0 = 1.093268816632711E-6
+ wa0 = 1.035196487524024E-5 pa0 = -4.928943147837386E-12 ags = -1.191493483525002
+ lags = 1.16248294127166E-6 wags = 1.21439877783786E-5 pags = -5.78218976484607E-12
+ b0 = 0 b1 = 0 keta = -0.081102291173502
+ lketa = 2.005927328052309E-8 wketa = -1.416725564926262E-7 pketa = 1.07605112780992E-13
+ a1 = 0 a2 = 0.42385546 rdsw = 65.968
+ rdswmin = 0 rdw = 0 rdwmin = 0
+ rsw = 0 rswmin = 0 prwb = 0
+ prwg = 0.021507 wr = 1 voff = -0.107048356364469
+ lvoff = -6.533844984870948E-9 wvoff = -4.157563510517169E-9 pvoff = -4.275527082103648E-14
+ voffl = 5.8197729E-9 minv = 0 nfactor = 2.540704899373772
+ lnfactor = 2.069684632785476E-7 wnfactor = -3.835168691235889E-7 pnfactor = -3.919759284290669E-13
+ eta0 = -0.451815060387666 leta0 = 4.484320555927418E-7 weta0 = -6.856480995916697E-8
+ peta0 = 3.264617435471792E-14 etab = 2.38360893990171E-4 letab = -2.622847026209041E-10
+ wetab = -3.831943721367735E-9 petab = 1.824526355717148E-15 dsub = -1.70710363277456
+ ldsub = 1.047052630861483E-6 wdsub = 1.27861286565513E-5 pdsub = -6.407414733876143E-12
+ cit = 0 cdsc = 0 cdscb = 0
+ cdscd = 5.4E-3 pclm = 0.265060463878963 lpclm = 2.623034990707567E-7
+ wpclm = -7.91883812691416E-8 ppclm = -8.875767192532802E-13 pdiblc1 = 0.679242722746118
+ lpdiblc1 = 2.961014292620497E-7 wpdiblc1 = -1.745617575554019E-6 ppdiblc1 = -1.662218554918302E-13
+ pdiblc2 = -1.452074581594853E-3 lpdiblc2 = 2.821978282547936E-9 wpdiblc2 = 4.188817167786844E-8
+ ppdiblc2 = -2.342040628954801E-14 pdiblcb = 0.022974484260031 lpdiblcb = -2.284237903763403E-8
+ wpdiblcb = 3.187895079876586E-9 ppdiblcb = -1.517871611752118E-15 drout = 1.020293090799388
+ ldrout = -7.421494564805513E-7 wdrout = -6.870374050996677E-6 pdrout = 6.706419444643692E-12
+ pscbe1 = -1.461636461476959E9 lpscbe1 = 680.7484247078605 wpscbe1 = 9.998067113033081E3
+ ppscbe1 = -2.797265732688057E-3 pscbe2 = 1E-12 pvag = 0
+ delta = 0.01 fprout = 0 pdits = 0
+ pditsl = 0 pditsd = 0 lambda = 0
+ vtl = 0 lc = 5E-9 xn = 3
+ alpha0 = -2.045363005314385E-5 lalpha0 = 1.963972049374442E-11 walpha0 = 1.383882472090581E-10
+ palpha0 = -1.14893032624048E-16 alpha1 = 0.916377248 lalpha1 = -3.160459735372802E-8
+ beta0 = 1.569617265101627 lbeta0 = 1.403287030115302E-5 wbeta0 = 9.041675895826209E-5
+ pbeta0 = -8.359790114360646E-11 aigbacc = 1 bigbacc = 0
+ cigbacc = 0 nigbacc = 0 aigbinv = 0.35
+ bigbinv = 0.03 cigbinv = 6E-3 eigbinv = 1.1
+ nigbinv = 0 aigc = 0.43 bigc = 0.054
+ cigc = 0.075 aigsd = 0.43 bigsd = 0.054
+ cigsd = 0.075 dlcig = 0 nigc = 0
+ poxedge = 1 pigcd = 1 ntox = 1
+ toxref = 4.148E-9 agidl = 0 bgidl = 2.3E9
+ cgidl = 0.5 egidl = 0.8 noia = 2.5E42
+ noib = 0 noic = 0 em = 4.1E7
+ af = 1 ef = 0.84 kf = 0
+ lintnoi = -1E-7 tnoia = 1.5E7 tnoib = 9.9E6
+ ntnoi = 1 rnoia = 0.94 rnoib = 0.26
+ xpart = 0 cgso = {2.449068E-10/sw_func_tox_lv_ratio} cgdo = {2.449068E-10/sw_func_tox_lv_ratio}
+ cgbo = {1E-13/sw_func_tox_lv_ratio} ckappas = 0.6 cf = 1.4067E-12
+ clc = 1E-7 cle = 0.6 dlc = 9.87908E-9
+ dwc = 0 vfbcv = -1 noff = 3.4037
+ voffcv = -0.17287 acde = 0.4 moin = 6.9
+ cgsl = {0/sw_func_tox_lv_ratio} cgdl = {0/sw_func_tox_lv_ratio} ijthsrev = 0.1
+ ijthsfwd = 0.1 xjbvs = 1 bvs = 11.7
+ jss = 2.75E-3 jsws = 6E-10 cjs = {sw_nsd_pw_cj}
+ mjs = 0.44 mjsws = 9E-4 cjsws = {3.67354204E-11*sw_func_nsd_pw_cj}
+ cjswgs = {2.38232788E-10*sw_func_nsd_pw_cj} mjswgs = 0.8 pbs = 0.729
+ pbsws = 0.2 pbswgs = 0.95578 xrcrg1 = 12
+ xrcrg2 = 1 rbpb = 50 rbpd = 50
+ rbps = 50 rbdb = 50 rbsb = 50
+ gbmin = 1E-12 tnom = 30 ute = -0.680326432762263
+ lute = -3.028715436078531E-7 wute = 2.142545093521423E-6 pute = -1.386698813274027E-12
+ kt1 = -0.268655366752023 lkt1 = -1.777383128919181E-9 wkt1 = -1.171499994328383E-9
+ pkt1 = -1.388875691723358E-14 kt1l = 0 kt2 = -0.017576666853973
+ lkt2 = -8.506170576148047E-9 wkt2 = 2.911051177726006E-9 pkt2 = -3.49345325361701E-15
+ ua1 = 2.58225373505154E-9 lua1 = -5.891710655620661E-16 wua1 = 4.53472896993511E-15
+ pua1 = -2.895121747011377E-21 ub1 = -1.239485764905863E-18 lub1 = -5.456547925937168E-26
+ wub1 = -3.366333664844644E-24 pub1 = 2.115558900144282E-30 uc1 = 1.498316505102567E-10
+ luc1 = -7.900978524043387E-17 wuc1 = -1.926657219579703E-16 puc1 = 9.963794597002815E-23
+ at = 7.989657715863558E4 lat = -0.013091084804129 wat = -0.049159335510696
+ pat = 2.680427210093172E-8 prt = 0 njs = 1.2928
+ xtis = 2 tpb = 1.2287E-3 tpbsw = 0
+ tpbswg = 0 tcj = 7.92E-4 tcjsw = 1E-5
+ tcjswg = 0 tvoff = 0 tvfbsdoff = 0
+ saref = 2.75E-6 sbref = 2.74E-6 wlod = 0
+ ku0 = -2.7E-8 kvsat = 0.2 kvth0 = 9.8E-9
+ tku0 = 0 llodku0 = 0 wlodku0 = 1
+ llodvth = 0 wlodvth = 1 lku0 = 0
+ wku0 = 0 pku0 = 0 lkvth0 = 0
+ wkvth0 = 2E-7 pkvth0 = 0 stk2 = 0
+ lodk2 = 1 steta0 = 0 lodeta0 = 1

.model nshort_model.14 nmos
+ level = 54 lmin = 2.5E-7 lmax = 5E-7 wmin = 5E-6
+ wmax = 7E-6 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 4.148E-9
+ toxm = 4.148E-9 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 9.999999999999999E22 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {2.1859E-8+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {1.1932E-8-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = 0 dwb = 0 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = 0.600055913168463 lvth0 = -1.836187806307696E-8
+ wvth0 = 1.376410745899428E-7 pvth0 = -1.834275596200204E-14 k1 = 0.282287833441199
+ lk1 = 1.065012081093659E-7 wk1 = -3.214225439102723E-7 pk1 = 8.60635555438369E-14
+ k2 = 0.052085107878465 lk2 = -3.093679873919933E-8 wk2 = 6.958429471233679E-8
+ pk2 = -1.897283581757019E-14 k3 = 2 k3b = 0.54
+ w0 = 0 lpe0 = 1.0325E-7 lpeb = -7.082E-8
+ vbm = -3 dvtp0 = 0 dvtp1 = 0
+ dvt0 = 0 dvt1 = 0.53 dvt2 = -0.032
+ dvt0w = -3.58 dvt1w = 1.6706E6 dvt2w = 0.068
+ vfbsdoff = 0 u0 = 0.026153897181042 lu0 = -1.70196903439523E-9
+ wu0 = 2.062968543927908E-8 pu0 = -6.263490726903066E-15 ua = -1.349419497710931E-9
+ lua = -1.867602033897232E-16 wua = 1.518287227989931E-15 pua = -2.777543678787653E-22
+ ub = 1.999102462218046E-18 lub = 1.765513674564946E-25 wub = -2.100701032220624E-25
+ pub = -2.383914575805439E-31 uc = 4.031218940556071E-12 luc = 3.891280702433506E-17
+ wuc = 5.360116115393456E-16 puc = -2.651788647166569E-22 ud = 0
+ up = 0 lp = 1 eu = 1.67
+ vsat = 4.89286190200102E4 lvsat = 0.021755806808461 wvsat = 0.299777690254014
+ pvsat = -7.952395718617654E-8 a0 = 1.5 ags = 2.363013911532893
+ lags = -5.299459917816256E-7 pags = 1.856110884906599E-18 b0 = 0
+ b1 = 0 keta = -0.025409731317712 lketa = -6.457959398973355E-9
+ wketa = 6.363471476463599E-8 pketa = 9.850929873644291E-15 a1 = 0
+ a2 = 0.42385546 rdsw = 65.968 rdswmin = 0
+ rdw = 0 rdwmin = 0 rsw = 0
+ rswmin = 0 prwb = 0 prwg = 0.021507
+ wr = 1 voff = -0.103106212294419 lvoff = -8.410841693808342E-9
+ wvoff = -1.66156889669133E-7 pvoff = 3.43784403388222E-14 voffl = 5.8197729E-9
+ minv = 0 nfactor = 3.336221670863461 lnfactor = -1.718057102314666E-7
+ wnfactor = -3.857714841000195E-6 pnfactor = 1.262214797108372E-12 eta0 = 0.49
+ etab = -2.569930338292707E-4 letab = -2.642886484466635E-11 wetab = 3.24661150286241E-9
+ petab = -1.545828614526896E-15 dsub = 0.387328261998424 ldsub = 4.981820621185383E-8
+ wdsub = -9.651936127768832E-7 pdsub = 1.400848461527026E-13 cit = 0
+ cdsc = 0 cdscb = 0 cdscd = 5.4E-3
+ pclm = 1.211362671563701 lpclm = -1.882650488874239E-7 wpclm = -3.909760515921197E-6
+ ppclm = 9.362965746514104E-13 pdiblc1 = 3.226103048537282 lpdiblc1 = -9.165504588188516E-7
+ wpdiblc1 = -9.936612420671622E-6 ppdiblc1 = 3.733805666083084E-12 pdiblc2 = 6.207590322382611E-3
+ lpdiblc2 = -8.250639261722778E-10 wpdiblc2 = -1.378271132350408E-8 ppdiblc2 = 3.086505259193493E-15
+ pdiblcb = 0.6042263145408 lpdiblcb = -2.995973005001984E-7 wpdiblcb = -3.118623056684907E-6
+ ppdiblcb = 1.484888707717725E-12 drout = -1.929948741598776 ldrout = 6.625668886301808E-7
+ wdrout = 1.374074810199336E-5 pdrout = -3.107277812792369E-12 pscbe1 = -7.843924540557315E8
+ lpscbe1 = 358.28817199034694 wpscbe1 = 7.852695800972251E3 ppscbe1 = -1.775777217648661E-3
+ pscbe2 = 1E-12 pvag = 0 delta = 0.01
+ fprout = 0 pdits = 0 pditsl = 0
+ pditsd = 0 lambda = 0 vtl = 0
+ lc = 5E-9 xn = 3 alpha0 = 4.138540030427234E-5
+ lalpha0 = -9.80406806451429E-12 walpha0 = -2.250088190308333E-10 palpha0 = 5.813339290714892E-17
+ alpha1 = 0.85 beta0 = 42.44059301879679 lbeta0 = -5.427272610308384E-6
+ wbeta0 = -1.665082017345302E-4 pbeta0 = 3.873332194081686E-11 aigbacc = 1
+ bigbacc = 0 cigbacc = 0 nigbacc = 0
+ aigbinv = 0.35 bigbinv = 0.03 cigbinv = 6E-3
+ eigbinv = 1.1 nigbinv = 0 aigc = 0.43
+ bigc = 0.054 cigc = 0.075 aigsd = 0.43
+ bigsd = 0.054 cigsd = 0.075 dlcig = 0
+ nigc = 0 poxedge = 1 pigcd = 1
+ ntox = 1 toxref = 4.148E-9 agidl = 0
+ bgidl = 2.3E9 cgidl = 0.5 egidl = 0.8
+ noia = 2.5E42 noib = 0 noic = 0
+ em = 4.1E7 af = 1 ef = 0.84
+ kf = 0 lintnoi = -1E-7 tnoia = 1.5E7
+ tnoib = 9.9E6 ntnoi = 1 rnoia = 0.94
+ rnoib = 0.26 xpart = 0 cgso = {2.449068E-10/sw_func_tox_lv_ratio}
+ cgdo = {2.449068E-10/sw_func_tox_lv_ratio} cgbo = {1E-13/sw_func_tox_lv_ratio} ckappas = 0.6
+ cf = 1.4067E-12 clc = 1E-7 cle = 0.6
+ dlc = 9.87908E-9 dwc = 0 vfbcv = -1
+ noff = 3.4037 voffcv = -0.17287 acde = 0.4
+ moin = 6.9 cgsl = {0/sw_func_tox_lv_ratio} cgdl = {0/sw_func_tox_lv_ratio}
+ ijthsrev = 0.1 ijthsfwd = 0.1 xjbvs = 1
+ bvs = 11.7 jss = 2.75E-3 jsws = 6E-10
+ cjs = {sw_nsd_pw_cj} mjs = 0.44 mjsws = 9E-4
+ cjsws = {3.67354204E-11*sw_func_nsd_pw_cj} cjswgs = {2.38232788E-10*sw_func_nsd_pw_cj} mjswgs = 0.8
+ pbs = 0.729 pbsws = 0.2 pbswgs = 0.95578
+ xrcrg1 = 12 xrcrg2 = 1 rbpb = 50
+ rbpd = 50 rbps = 50 rbdb = 50
+ rbsb = 50 gbmin = 1E-12 tnom = 30
+ ute = -1.212504930609545 lute = -4.948220235683988E-8 wute = -5.005194258228292E-6
+ pute = 2.016597210710675E-12 kt1 = -0.214382781580876 lkt1 = -2.761851474196813E-8
+ wkt1 = -3.400134791641692E-7 pkt1 = 1.474461076767777E-13 kt1l = 0
+ kt2 = -1.06813707072801E-3 lkt2 = -1.636647591302327E-8 wkt2 = -2.191664868057459E-7
+ pkt2 = 1.022456573716814E-13 ua1 = 1.746611269392912E-9 lua1 = -1.912916045332303E-16
+ wua1 = -6.466229626036761E-15 pua1 = 2.342830675040287E-21 ub1 = -2.10365655267725E-18
+ lub1 = 3.568973429469456E-25 wub1 = 3.572949935601235E-24 pub1 = -1.188483836237617E-30
+ uc1 = -1.358491247538446E-10 luc1 = 5.701311637071426E-17 wuc1 = 1.96502115319418E-16
+ puc1 = -8.565887139987843E-23 at = 7.917893228981526E4 lat = -0.012749388246868
+ wat = -6.070965093290702E-3 pat = 6.288347763870249E-9 prt = 0
+ njs = 1.2928 xtis = 2 tpb = 1.2287E-3
+ tpbsw = 0 tpbswg = 0 tcj = 7.92E-4
+ tcjsw = 1E-5 tcjswg = 0 tvoff = 0
+ tvfbsdoff = 0 saref = 1.75E-6 sbref = 1.74E-6
+ wlod = 0 ku0 = -2.7E-8 kvsat = 0.2
+ kvth0 = 9.8E-9 tku0 = 0 llodku0 = 0
+ wlodku0 = 1 llodvth = 0 wlodvth = 1
+ lku0 = 0 wku0 = 0 pku0 = 0
+ lkvth0 = 0 wkvth0 = 2E-7 pkvth0 = 0
+ stk2 = 0 lodk2 = 1 steta0 = 0
+ lodeta0 = 1

.model nshort_model.15 nmos
+ level = 54 lmin = 1.8E-7 lmax = 2.5E-7 wmin = 5E-6
+ wmax = 7E-6 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 4.148E-9
+ toxm = 4.148E-9 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 9.999999999999999E22 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {2.1859E-8+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {1.1932E-8-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = 0 dwb = 0 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = 0.586049365553648 lvth0 = -1.519449341165325E-8
+ wvth0 = 4.902589364002621E-7 pvth0 = -9.808234876034039E-14 k1 = 0.458080632459477
+ lk1 = 6.674812771056861E-8 wk1 = 1.733198695920878E-7 pk1 = -2.581551487593278E-14
+ k2 = 0.015994475136665 lk2 = -2.277540741349972E-8 wk2 = -1.488644617488886E-7
+ pk2 = 3.042629217354547E-14 k3 = 2 k3b = 0.54
+ w0 = 0 lpe0 = 1.0325E-7 lpeb = -7.082E-8
+ vbm = -3 dvtp0 = 0 dvtp1 = 0
+ dvt0 = 0 dvt1 = 0.53 dvt2 = -0.032
+ dvt0w = -3.58 dvt1w = 1.6706E6 dvt2w = 0.068
+ vfbsdoff = 0 u0 = -0.013794402535433 lu0 = 7.331779670289558E-9
+ wu0 = 3.161274109522536E-8 pu0 = -8.747155000716134E-15 ua = -5.194822301130732E-9
+ lua = 6.828238049644167E-16 wua = 8.593040434012419E-17 pua = 4.61530747941074E-23
+ ub = 4.384694129626147E-18 lub = -3.629167898445035E-25 wub = 2.765827802869489E-24
+ pub = -9.113491064724628E-31 uc = 3.482642912074568E-10 luc = -3.893068300581279E-17
+ wuc = -1.862306270780954E-15 puc = 2.771671479197262E-22 ud = 0
+ up = 0 lp = 1 eu = 1.67
+ vsat = 6.842631279793417E4 lvsat = 0.017346676328297 wvsat = 0.319214473473154
+ pvsat = -8.391931359622011E-8 a0 = 1.5 ags = -2.725049684046048
+ lags = 6.206483574682137E-7 wags = 1.39224243602144E-11 pags = -2.173791649906436E-18
+ b0 = 0 b1 = 0 keta = -0.113230348385952
+ lketa = 1.340144366237034E-8 wketa = 5.300964428252111E-7 pketa = -9.563285946306191E-14
+ a1 = 0 a2 = 0.42385546 rdsw = 65.968
+ rdswmin = 0 rdw = 0 rdwmin = 0
+ rsw = 0 rswmin = 0 prwb = 0
+ prwg = 0.021507 wr = 1 voff = -0.060728984567992
+ lvoff = -1.799385846295151E-8 wvoff = -3.732545738501178E-7 pvoff = 8.121068224877339E-14
+ voffl = 5.8197729E-9 minv = 0 nfactor = 2.261485731631155
+ lnfactor = 7.12307761227699E-8 wnfactor = -1.371177435903804E-6 pnfactor = 6.999191744694951E-13
+ eta0 = 1.550355063229624 leta0 = -2.397844525784943E-7 weta0 = -2.539778354749154E-7
+ peta0 = 5.743353180295545E-14 etab = 0.079519448489995 letab = -1.806675424527615E-8
+ wetab = -1.331586887207779E-7 petab = 2.930032035684622E-14 dsub = 1.052696561220498
+ ldsub = -1.006455195010292E-7 wdsub = -9.748341775119966E-7 pdsub = 1.422649248996422E-13
+ cit = 0 cdsc = 0 cdscb = 0
+ cdscd = 8.522720000000001E-3 lcdscd = -7.061594099200002E-10 pclm = 1.175664524230347
+ lpclm = -1.801924126420486E-7 wpclm = -3.364135541334164E-6 ppclm = 8.129111253981976E-13
+ pdiblc1 = -3.504829722811056 lpdiblc1 = 6.05555754362776E-7 wpdiblc1 = 2.12192708358484E-5
+ ppdiblc1 = -3.311661150013328E-12 pdiblc2 = -8.867346783530187E-3 lpdiblc2 = 2.583922051210418E-9
+ wpdiblc2 = -1.823973297898594E-8 ppdiblc2 = 4.09439830827754E-15 pdiblcb = -2.245021455576421
+ lpdiblcb = 3.447201932430297E-7 wpdiblcb = 1.190062844236073E-5 ppdiblcb = -1.911504749270459E-12
+ drout = 2.107148648874746 ldrout = -2.503661668619396E-7 wdrout = -3.309056972963674E-6
+ pdrout = 7.482969076381133E-13 pscbe1 = 8.184696981923373E8 lpscbe1 = -4.176663670422391
+ wpscbe1 = -64.81001347413296 ppscbe1 = 1.465587720698653E-5 pscbe2 = 1E-12
+ pvag = 0 delta = 0.01 fprout = 0
+ pdits = 0 pditsl = 0 pditsd = 0
+ lambda = 0 vtl = 0 lc = 5E-9
+ xn = 3 alpha0 = 3.095849207334765E-6 lalpha0 = -1.145422137657215E-12
+ walpha0 = 3.763936371948774E-11 palpha0 = -1.260816547277671E-18 alpha1 = -2.783651019360897
+ lalpha1 = 8.216993069141955E-7 walpha1 = 1.998416411725231E-5 palpha1 = -4.519138936818969E-12
+ beta0 = 44.86413993147485 lbeta0 = -5.975323814953751E-6 wbeta0 = -1.149999147611612E-4
+ pbeta0 = 2.708544395780709E-11 aigbacc = 1 bigbacc = 0
+ cigbacc = 0 nigbacc = 0 aigbinv = 0.35
+ bigbinv = 0.03 cigbinv = 6E-3 eigbinv = 1.1
+ nigbinv = 0 aigc = 0.43 bigc = 0.054
+ cigc = 0.075 aigsd = 0.43 bigsd = 0.054
+ cigsd = 0.075 dlcig = 0 nigc = 0
+ poxedge = 1 pigcd = 1 ntox = 1
+ toxref = 4.148E-9 agidl = 0 bgidl = 2.3E9
+ cgidl = 0.5 egidl = 0.8 noia = 2.5E42
+ noib = 0 noic = 0 em = 4.1E7
+ af = 1 ef = 0.84 kf = 0
+ lintnoi = -1E-7 tnoia = 1.5E7 tnoib = 9.9E6
+ ntnoi = 1 rnoia = 0.94 rnoib = 0.26
+ xpart = 0 cgso = {2.449068E-10/sw_func_tox_lv_ratio} cgdo = {2.449068E-10/sw_func_tox_lv_ratio}
+ cgbo = {1E-13/sw_func_tox_lv_ratio} ckappas = 0.6 cf = 1.4067E-12
+ clc = 1E-7 cle = 0.6 dlc = 9.87908E-9
+ dwc = 0 vfbcv = -1 noff = 3.4037
+ voffcv = -0.17287 acde = 0.4 moin = 6.9
+ cgsl = {0/sw_func_tox_lv_ratio} cgdl = {0/sw_func_tox_lv_ratio} ijthsrev = 0.1
+ ijthsfwd = 0.1 xjbvs = 1 bvs = 11.7
+ jss = 2.75E-3 jsws = 6E-10 cjs = {sw_nsd_pw_cj}
+ mjs = 0.44 mjsws = 9E-4 cjsws = {3.67354204E-11*sw_func_nsd_pw_cj}
+ cjswgs = {2.38232788E-10*sw_func_nsd_pw_cj} mjswgs = 0.8 pbs = 0.729
+ pbsws = 0.2 pbswgs = 0.95578 xrcrg1 = 12
+ xrcrg2 = 1 rbpb = 50 rbpd = 50
+ rbps = 50 rbdb = 50 rbsb = 50
+ gbmin = 1E-12 tnom = 30 ute = -0.605933312298173
+ lute = -1.866498818353003E-7 wute = 1.299739769783044E-5 pute = -2.054436923864622E-12
+ kt1 = -0.584844743242046 lkt1 = 5.615627142024206E-8 wkt1 = 1.534668965145515E-6
+ pkt1 = -2.764870815496369E-13 kt1l = 0 kt2 = -0.155359043103535
+ lkt2 = 1.852425241361149E-8 wkt2 = 7.440012127551652E-7 pkt2 = -1.155612335362248E-13
+ ua1 = 4.223758656352509E-9 lua1 = -7.514638060307257E-16 wua1 = 1.204986546830962E-14
+ pua1 = -1.844325005214825E-21 ub1 = -4.489634735145902E-18 lub1 = 8.964529052176764E-25
+ wub1 = -2.407922044394457E-25 pub1 = -3.260594436573779E-31 uc1 = -9.851794355482102E-11
+ luc1 = 4.857119237909186E-17 wuc1 = 6.668615294827137E-16 puc1 = -1.920240678811094E-22
+ at = 3.846530240548508E4 lat = -3.54257083934544E-3 wat = -0.24305069202783
+ pat = 5.987799529393932E-8 prt = 0 njs = 1.2928
+ xtis = 2 tpb = 1.2287E-3 tpbsw = 0
+ tpbswg = 0 tcj = 7.92E-4 tcjsw = 1E-5
+ tcjswg = 0 tvoff = 0 tvfbsdoff = 0
+ saref = 1.25E-6 sbref = 1.24E-6 wlod = 0
+ ku0 = -2.7E-8 kvsat = 0.2 kvth0 = 9.8E-9
+ tku0 = 0 llodku0 = 0 wlodku0 = 1
+ llodvth = 0 wlodvth = 1 lku0 = 0
+ wku0 = 0 pku0 = 0 lkvth0 = 0
+ wkvth0 = 2E-7 pkvth0 = 0 stk2 = 0
+ lodk2 = 1 steta0 = 0 lodeta0 = 1

.model nshort_model.16 nmos
+ level = 54 lmin = 1.5E-7 lmax = 1.8E-7 wmin = 5E-6
+ wmax = 7E-6 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 4.148E-9
+ toxm = 4.148E-9 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 9.999999999999999E22 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {2.1859E-8+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {1.1932E-8-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = 0 dwb = 0 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = 0.497680789006495 lvth0 = -1.396977343886954E-9
+ wvth0 = 6.757248245883855E-7 pvth0 = -1.270402506784811E-13 k1 = 0.80245941064215
+ lk1 = 1.297820280023876E-8 wk1 = 1.181647507247276E-7 pk1 = -1.720381523645863E-14
+ k2 = -0.022428797958142 lk2 = -1.6776151245569E-8 wk2 = -4.839081426772983E-7
+ pk2 = 8.273867233898364E-14 k3 = 2 k3b = 0.54
+ w0 = 0 lpe0 = 1.0325E-7 lpeb = -7.082E-8
+ vbm = -3 dvtp0 = 0 dvtp1 = 0
+ dvt0 = 0 dvt1 = 0.53 dvt2 = -0.032
+ dvt0w = -3.58 dvt1w = 1.6706E6 dvt2w = 0.068
+ vfbsdoff = 0 u0 = 0.068621224186513 lu0 = -5.536266623568184E-9
+ wu0 = 9.414146324922376E-8 pu0 = -1.851013956295283E-14 ua = 6.033562109762451E-9
+ lua = -1.070331223414801E-15 wua = 4.584847861296159E-16 pua = -1.201607616097668E-23
+ ub = -5.14963473875173E-18 lub = 1.125735182348545E-24 wub = 6.867891660182195E-24
+ pub = -1.551828948897839E-30 uc = 1.721098632245748E-10 luc = -1.142663523827753E-17
+ wuc = 3.768785961303405E-16 puc = -7.245022046033562E-23 ud = 0
+ up = 0 lp = 1 eu = 1.67
+ vsat = 2.279489769160281E5 lvsat = -7.560554356445911E-3 wvsat = -1.046666644325516
+ pvsat = 1.29343900612393E-7 a0 = 1.5 ags = 1.25
+ b0 = 0 b1 = 0 keta = -1.086656882003298
+ lketa = 1.653883689152482E-7 wketa = 5.4800403457398E-6 pketa = -8.68497300688534E-13
+ a1 = 0 a2 = 0.42385546 rdsw = 65.968
+ rdswmin = 0 rdw = 0 rdwmin = 0
+ rsw = 0 rswmin = 0 prwb = 0
+ prwg = 0.021507 wr = 1 voff = 0.55466020051224
+ lvoff = -1.140782642646386E-7 wvoff = -3.093003668120484E-6 pvoff = 5.058614268317713E-13
+ voffl = 5.8197729E-9 minv = 0 nfactor = 28.041128670414697
+ lnfactor = -3.953899553767136E-6 wnfactor = -1.224818552693739E-4 pnfactor = 1.960965596867618E-11
+ eta0 = 0.072061156477103 leta0 = -8.969555153782614E-9 weta0 = 5.975626640990564E-7
+ peta0 = -7.552259563852616E-14 etab = 0.03506506218337 letab = -1.112582418490492E-8
+ wetab = -2.497332409541006E-8 petab = 1.240869026569979E-14 dsub = 1.43959292470115
+ ldsub = -1.610539701094443E-7 wdsub = -5.121179047785371E-6 pdsub = 7.896586275646457E-13
+ cit = 0 cdsc = 0 cdscb = 0
+ cdscd = 0.027579751562142 lcdscd = -3.681648089906581E-9 wcdscd = -1.05531562266066E-7
+ pcdscd = 1.647727600597448E-14 pclm = -0.871159991646503 lpclm = 1.393905799688993E-7
+ wpclm = 1.147277413387082E-5 ppclm = -1.503664603649607E-12 pdiblc1 = -0.128069597134514
+ lpdiblc1 = 7.832193538014348E-8 wpdiblc1 = 3.15245767976486E-6 ppdiblc1 = -4.907812110750675E-13
+ pdiblc2 = -6.906294731612566E-3 lpdiblc2 = 2.277731228032208E-9 wpdiblc2 = 8.833404804172024E-8
+ ppdiblc2 = -1.254560556517144E-14 pdiblcb = -0.56672302415965 lpdiblcb = 8.267738935534055E-8
+ wpdiblcb = 8.161113284529011E-7 ppdiblcb = -1.808125851733463E-13 drout = -0.248743257952596
+ ldrout = 1.174733719024542E-7 wdrout = 1.199121754639496E-5 pdrout = -1.640626754716466E-12
+ pscbe1 = 8.143741680702468E8 lpscbe1 = -3.537203979279664 wpscbe1 = 28.25952500649075
+ ppscbe1 = 1.243717467758651E-7 pscbe2 = 1E-12 pvag = 0
+ delta = 0.01 fprout = 0 pdits = 0
+ pditsl = 0 pditsd = 0 lambda = 0
+ vtl = 0 lc = 5E-9 xn = 3
+ alpha0 = -2.219442352735979E-5 lalpha0 = 2.803299886047054E-12 walpha0 = 1.538681048809421E-10
+ palpha0 = -1.940830727726251E-17 alpha1 = 9.328519045175417 lalpha1 = -1.069446478282246E-6
+ walpha1 = -4.66297162735887E-5 palpha1 = 5.881685891885382E-12 beta0 = -23.95538075376639
+ lbeta0 = 4.769880866757076E-6 wbeta0 = 3.043272422219475E-4 pbeta0 = -3.838662102490757E-11
+ aigbacc = 1 bigbacc = 0 cigbacc = 0
+ nigbacc = 0 aigbinv = 0.35 bigbinv = 0.03
+ cigbinv = 6E-3 eigbinv = 1.1 nigbinv = 0
+ aigc = 0.43 bigc = 0.054 cigc = 0.075
+ aigsd = 0.43 bigsd = 0.054 cigsd = 0.075
+ dlcig = 0 nigc = 0 poxedge = 1
+ pigcd = 1 ntox = 1 toxref = 4.148E-9
+ agidl = 0 bgidl = 2.3E9 cgidl = 0.5
+ egidl = 0.8 noia = 2.5E42 noib = 0
+ noic = 0 em = 4.1E7 af = 1
+ ef = 0.84 kf = 0 lintnoi = -1E-7
+ tnoia = 1.5E7 tnoib = 9.9E6 ntnoi = 1
+ rnoia = 0.94 rnoib = 0.26 xpart = 0
+ cgso = {2.449068E-10/sw_func_tox_lv_ratio} cgdo = {2.449068E-10/sw_func_tox_lv_ratio} cgbo = {1E-13/sw_func_tox_lv_ratio}
+ ckappas = 0.6 cf = 1.4067E-12 clc = 1E-7
+ cle = 0.6 dlc = 9.87908E-9 dwc = 0
+ vfbcv = -1 noff = 3.4037 voffcv = -0.17287
+ acde = 0.4 moin = 6.9 cgsl = {0/sw_func_tox_lv_ratio}
+ cgdl = {0/sw_func_tox_lv_ratio} ijthsrev = 0.1 ijthsfwd = 0.1
+ xjbvs = 1 bvs = 11.7 jss = 2.75E-3
+ jsws = 6E-10 cjs = {sw_nsd_pw_cj} mjs = 0.44
+ mjsws = 9E-4 cjsws = {3.67354204E-11*sw_func_nsd_pw_cj} cjswgs = {2.38232788E-10*sw_func_nsd_pw_cj}
+ mjswgs = 0.8 pbs = 0.729 pbsws = 0.2
+ pbswgs = 0.95578 xrcrg1 = 12 xrcrg2 = 1
+ rbpb = 50 rbpd = 50 rbps = 50
+ rbdb = 50 rbsb = 50 gbmin = 1E-12
+ tnom = 30 ute = -9.375262849476252 lute = 1.182558154781536E-6
+ wute = -8.358412305389467E-7 pute = 1.054296694552606E-13 kt1 = -0.526935792087742
+ lkt1 = 4.71145994228138E-8 wkt1 = 5.845589058150978E-7 pkt1 = -1.281406973260229E-13
+ kt1l = 0 kt2 = -0.064724877300995 lkt2 = 4.372996301866103E-9
+ wkt2 = 1.930320397133724E-9 pkt2 = 3.02747312988792E-16 ua1 = -1.32110960650442E-8
+ lua1 = 1.970744670749271E-15 wua1 = 1.372150594674625E-14 pua1 = -2.105328262956007E-21
+ ub1 = 8.031610842555904E-18 lub1 = -1.058564294302372E-24 wub1 = -6.900660489851569E-24
+ pub1 = 7.137857509537293E-31 uc1 = 2.439604407897182E-10 luc1 = -4.90201263892711E-18
+ wuc1 = -1.576303213044202E-15 puc1 = 1.582147023580731E-22 at = 2.162270651606062E5
+ lat = -0.031297581428879 wat = -1.159255683299305 pat = 2.029305778111023E-7
+ prt = 0 njs = 1.2928 xtis = 2
+ tpb = 1.2287E-3 tpbsw = 0 tpbswg = 0
+ tcj = 7.92E-4 tcjsw = 1E-5 tcjswg = 0
+ tvoff = 0 tvfbsdoff = 0 saref = 1.1E-6
+ sbref = 1.1E-6 wlod = 0 ku0 = -2.7E-8
+ kvsat = 0.2 kvth0 = 9.8E-9 tku0 = 0
+ llodku0 = 0 wlodku0 = 1 llodvth = 0
+ wlodvth = 1 lku0 = 0 wku0 = 0
+ pku0 = 0 lkvth0 = 0 wkvth0 = 2E-7
+ pkvth0 = 0 stk2 = 0 lodk2 = 1
+ steta0 = 0 lodeta0 = 1

.model nshort_model.17 nmos
+ level = 54 lmin = 8E-6 lmax = 2.02E-5 wmin = 3E-6
+ wmax = 5E-6 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 4.148E-9
+ toxm = 4.148E-9 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 9.999999999999999E22 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {2.1859E-8+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {1.1932E-8-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = 0 dwb = 0 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = 0.5144028148889 wvth0 = 2.137091856221296E-8
+ k1 = 0.52900534172472 wk1 = 6.64042081249815E-8 k2 = -0.022170206002009
+ wk2 = -2.271709375563281E-8 k3 = 2 k3b = 0.54
+ w0 = 0 lpe0 = 1.0325E-7 lpeb = -7.082E-8
+ vbm = -3 dvtp0 = 0 dvtp1 = 0
+ dvt0 = 0 dvt1 = 0.53 dvt2 = -0.032
+ dvt0w = -3.58 dvt1w = 1.6706E6 dvt2w = 0.068
+ vfbsdoff = 0 u0 = 0.0321517281211 wu0 = -3.861578682301743E-9
+ ua = -7.486422007807401E-10 wua = 1.29680032017528E-16 ub = 1.65683489561E-18
+ wub = -3.385383246237228E-25 uc = 1.102824735099999E-11 wuc = 1.77210636968691E-16
+ ud = 0 up = 0 lp = 1
+ eu = 1.67 vsat = 8E4 a0 = 1.2646697222779
+ wa0 = 4.658517385848453E-7 ags = 0.3785123705454 wags = 1.082106508913035E-7
+ b0 = -3.114886529299998E-24 wb0 = 1.543825603721206E-29 b1 = 0
+ keta = -6.9689624785628E-3 wketa = 3.87587040625059E-9 a1 = 0
+ a2 = 0.42385546 rdsw = 65.968 rdswmin = 0
+ rdw = 0 rdwmin = 0 rsw = 0
+ rswmin = 0 prwb = 0 prwg = 0.021507
+ wr = 1 voff = -0.10161544947289 wvoff = -1.221778293352582E-8
+ voffl = 5.8197729E-9 minv = 0 nfactor = 2.71425
+ eta0 = 0.08 etab = -0.07 dsub = 0.56
+ cit = 0 cdsc = 0 cdscb = 0
+ cdscd = 5.4E-3 pclm = 0.067053840491 wpclm = 4.871113006758543E-8
+ pdiblc1 = 0.39 pdiblc2 = 4.2744340571756E-3 wpdiblc2 = -5.356477769096595E-9
+ pdiblcb = 3.650569947740599 wpdiblcb = -1.821716117172767E-5 drout = 0.56
+ pscbe1 = 5.482158036073201E8 wpscbe1 = 725.1759048101046 pscbe2 = 1E-12
+ pvag = 0 delta = 0.01 fprout = 0
+ pdits = 0 pditsl = 0 pditsd = 0
+ lambda = 0 vtl = 0 lc = 5E-9
+ xn = 3 alpha0 = 3E-8 alpha1 = 0.85
+ beta0 = 13.86 aigbacc = 1 bigbacc = 0
+ cigbacc = 0 nigbacc = 0 aigbinv = 0.35
+ bigbinv = 0.03 cigbinv = 6E-3 eigbinv = 1.1
+ nigbinv = 0 aigc = 0.43 bigc = 0.054
+ cigc = 0.075 aigsd = 0.43 bigsd = 0.054
+ cigsd = 0.075 dlcig = 0 nigc = 0
+ poxedge = 1 pigcd = 1 ntox = 1
+ toxref = 4.148E-9 agidl = 0 bgidl = 2.3E9
+ cgidl = 0.5 egidl = 0.8 noia = 2.5E42
+ noib = 0 noic = 0 em = 4.1E7
+ af = 1 ef = 0.84 kf = 0
+ lintnoi = -1E-7 tnoia = 1.5E7 tnoib = 9.9E6
+ ntnoi = 1 rnoia = 0.94 rnoib = 0.26
+ xpart = 0 cgso = {2.449068E-10/sw_func_tox_lv_ratio} cgdo = {2.449068E-10/sw_func_tox_lv_ratio}
+ cgbo = {1E-13/sw_func_tox_lv_ratio} ckappas = 0.6 cf = 1.4067E-12
+ clc = 1E-7 cle = 0.6 dlc = 9.87908E-9
+ dwc = 0 vfbcv = -1 noff = 3.4037
+ voffcv = -0.17287 acde = 0.4 moin = 6.9
+ cgsl = {0/sw_func_tox_lv_ratio} cgdl = {0/sw_func_tox_lv_ratio} ijthsrev = 0.1
+ ijthsfwd = 0.1 xjbvs = 1 bvs = 11.7
+ jss = 2.75E-3 jsws = 6E-10 cjs = {sw_nsd_pw_cj}
+ mjs = 0.44 mjsws = 9E-4 cjsws = {3.67354204E-11*sw_func_nsd_pw_cj}
+ cjswgs = {2.38232788E-10*sw_func_nsd_pw_cj} mjswgs = 0.8 pbs = 0.729
+ pbsws = 0.2 pbswgs = 0.95578 xrcrg1 = 12
+ xrcrg2 = 1 rbpb = 50 rbpd = 50
+ rbps = 50 rbdb = 50 rbsb = 50
+ gbmin = 1E-12 tnom = 30 ute = -2.0217583694
+ wute = 6.842562112065701E-7 kt1 = -0.33631381646 wkt1 = 5.904823407200179E-8
+ kt1l = 0 kt2 = -0.052084039143581 wkt2 = 3.258525514677992E-8
+ ua1 = 1.529990390200001E-10 wua1 = 5.258662830878761E-16 ub1 = -6.0529606929E-19
+ wub1 = 5.325330191927798E-25 uc1 = 1.977567061289501E-11 wuc1 = -1.362354849120647E-17
+ at = 1.4E5 prt = 0 njs = 1.2928
+ xtis = 2 tpb = 1.2287E-3 tpbsw = 0
+ tpbswg = 0 tcj = 7.92E-4 tcjsw = 1E-5
+ tcjswg = 0 tvoff = 0 tvfbsdoff = 0
+ saref = 3E-6 sbref = 3E-6 wlod = 0
+ ku0 = -2.7E-8 kvsat = 0.2 kvth0 = 9.8E-9
+ tku0 = 0 llodku0 = 0 wlodku0 = 1
+ llodvth = 0 wlodvth = 1 lku0 = 0
+ wku0 = 0 pku0 = 0 lkvth0 = 0
+ wkvth0 = 2E-7 pkvth0 = 0 stk2 = 0
+ lodk2 = 1 steta0 = 0 lodeta0 = 1

.model nshort_model.18 nmos
+ level = 54 lmin = 4E-6 lmax = 8E-6 wmin = 3E-6
+ wmax = 5E-6 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 4.148E-9
+ toxm = 4.148E-9 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 9.999999999999999E22 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {2.1859E-8+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {1.1932E-8-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = 0 dwb = 0 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = 0.509404849246972 lvth0 = 3.986445368334391E-8
+ wvth0 = 1.28214088836722E-8 pvth0 = 6.81920519293574E-14 k1 = 0.514358429772291
+ lk1 = 1.168257617126003E-7 wk1 = 1.004324218257689E-7 pk1 = -2.714136603145434E-13
+ k2 = -0.014808763207177 lk2 = -5.871586888779976E-8 wk2 = -3.298876160905455E-8
+ pk2 = 8.19282197457199E-14 k3 = 2 k3b = 0.54
+ w0 = 0 lpe0 = 1.0325E-7 lpeb = -7.082E-8
+ vbm = -3 dvtp0 = 0 dvtp1 = 0
+ dvt0 = 0 dvt1 = 0.53 dvt2 = -0.032
+ dvt0w = -3.58 dvt1w = 1.6706E6 dvt2w = 0.068
+ vfbsdoff = 0 u0 = 0.031635376905427 lu0 = 4.118487519975638E-9
+ wu0 = -1.896065341383374E-9 pu0 = -1.567720171697927E-14 ua = -6.610039312395343E-10
+ lua = -6.990147566653148E-16 wua = -2.620612687561674E-16 pua = 3.124581891787901E-21
+ ub = 1.468911820506135E-18 lub = 1.498900004566642E-24 wub = 4.223971662712666E-25
+ pub = -6.069324962605197E-30 uc = -1.023161189022321E-10 luc = 9.040500800695901E-16
+ wuc = 5.426329931522462E-16 puc = -2.914658410360478E-21 ud = 0
+ up = 0 lp = 1 eu = 1.67
+ vsat = 8E4 a0 = 1.014825383465242 la0 = 1.992792425199841E-6
+ wa0 = 1.617523853630661E-6 pa0 = -9.18589341701307E-12 ags = 0.229018537540286
+ lags = 1.192383143210082E-6 wags = 5.315752334439462E-7 pags = -3.376813488023105E-12
+ b0 = -6.211189645566194E-24 lb0 = 2.469653475256299E-29 wb0 = 3.078440743890611E-29
+ pb0 = -1.224029906565024E-34 b1 = 0 keta = -9.975873028045135E-3
+ lketa = 2.398352748250585E-8 wketa = -1.84450310991871E-9 pketa = 4.562647713576453E-14
+ a1 = 0 a2 = 0.42385546 rdsw = 65.968
+ rdswmin = 0 rdw = 0 rdwmin = 0
+ rsw = 0 rswmin = 0 prwb = 0
+ prwg = 0.021507 wr = 1 voff = -0.101696598611351
+ lvoff = 6.472565646451855E-10 wvoff = -1.79817108853726E-8 pvoff = 4.59738732381313E-14
+ voffl = 5.8197729E-9 minv = 0 nfactor = 2.90364279197379
+ lnfactor = -1.54382952880319E-6 wnfactor = -7.580219357133228E-7 pnfactor = 6.144254900415152E-12
+ eta0 = 0.08 etab = -0.07 dsub = 0.56
+ cit = 0 cdsc = 0 cdscb = 0
+ cdscd = 5.4E-3 pclm = -0.355723849233697 lpclm = 3.372132351009984E-6
+ wpclm = 1.074726237610647E-7 ppclm = -4.686896652623327E-13 pdiblc1 = 0.39
+ pdiblc2 = 5.687552554288154E-3 lpdiblc2 = -1.127122531708533E-8 wpdiblc2 = -1.255694473117526E-8
+ ppdiblc2 = 5.743190375304623E-14 pdiblcb = 7.30421144517298 lpdiblcb = -2.914194147876432E-5
+ wpdiblcb = -3.632563875990482E-5 ppdiblcb = 1.444356799962529E-10 drout = 0.56
+ pscbe1 = 3.005663899936626E8 lpscbe1 = 1.975285403302784E3 wpscbe1 = 1.438242589061678E3
+ ppscbe1 = -5.687516850659606E-3 pscbe2 = 1E-12 pvag = 0
+ delta = 0.01 fprout = 0 pdits = 0
+ pditsl = 0 pditsd = 0 lambda = 0
+ vtl = 0 lc = 5E-9 xn = 3
+ alpha0 = 3E-8 alpha1 = 0.85 beta0 = 13.86
+ aigbacc = 1 bigbacc = 0 cigbacc = 0
+ nigbacc = 0 aigbinv = 0.35 bigbinv = 0.03
+ cigbinv = 6E-3 eigbinv = 1.1 nigbinv = 0
+ aigc = 0.43 bigc = 0.054 cigc = 0.075
+ aigsd = 0.43 bigsd = 0.054 cigsd = 0.075
+ dlcig = 0 nigc = 0 poxedge = 1
+ pigcd = 1 ntox = 1 toxref = 4.148E-9
+ agidl = 0 bgidl = 2.3E9 cgidl = 0.5
+ egidl = 0.8 noia = 2.5E42 noib = 0
+ noic = 0 em = 4.1E7 af = 1
+ ef = 0.84 kf = 0 lintnoi = -1E-7
+ tnoia = 1.5E7 tnoib = 9.9E6 ntnoi = 1
+ rnoia = 0.94 rnoib = 0.26 xpart = 0
+ cgso = {2.449068E-10/sw_func_tox_lv_ratio} cgdo = {2.449068E-10/sw_func_tox_lv_ratio} cgbo = {1E-13/sw_func_tox_lv_ratio}
+ ckappas = 0.6 cf = 1.4067E-12 clc = 1E-7
+ cle = 0.6 dlc = 9.87908E-9 dwc = 0
+ vfbcv = -1 noff = 3.4037 voffcv = -0.17287
+ acde = 0.4 moin = 6.9 cgsl = {0/sw_func_tox_lv_ratio}
+ cgdl = {0/sw_func_tox_lv_ratio} ijthsrev = 0.1 ijthsfwd = 0.1
+ xjbvs = 1 bvs = 11.7 jss = 2.75E-3
+ jsws = 6E-10 cjs = {sw_nsd_pw_cj} mjs = 0.44
+ mjsws = 9E-4 cjsws = {3.67354204E-11*sw_func_nsd_pw_cj} cjswgs = {2.38232788E-10*sw_func_nsd_pw_cj}
+ mjswgs = 0.8 pbs = 0.729 pbsws = 0.2
+ pbswgs = 0.95578 xrcrg1 = 12 xrcrg2 = 1
+ rbpb = 50 rbpd = 50 rbps = 50
+ rbdb = 50 rbsb = 50 gbmin = 1E-12
+ tnom = 30 ute = -2.363712446899473 lute = 2.727472227890337E-6
+ wute = 1.614943891715514E-6 pute = -7.42329151326389E-12 kt1 = -0.357459679754327
+ lkt1 = 1.68662281472962E-7 wkt1 = 1.280851606074074E-7 pkt1 = -5.506479150684042E-13
+ kt1l = 0 kt2 = -0.062500179452259 lkt2 = 8.308055169709611E-8
+ wkt2 = 6.661110935767231E-8 pkt2 = -2.713948407022504E-13 ua1 = -4.847675259755835E-10
+ lua1 = 5.086912858657615E-15 wua1 = 2.541307231229891E-15 pua1 = -1.607543110234966E-20
+ ub1 = -1.851937603054501E-19 lub1 = -3.350793150374793E-24 wub1 = -9.281076705424573E-25
+ pub1 = 1.165026878846206E-29 uc1 = 2.77605289039067E-11 luc1 = -6.36883156698369E-17
+ wuc1 = -7.244529656550389E-17 puc1 = 4.691702623983344E-22 at = 1.4E5
+ prt = 0 njs = 1.2928 xtis = 2
+ tpb = 1.2287E-3 tpbsw = 0 tpbswg = 0
+ tcj = 7.92E-4 tcjsw = 1E-5 tcjswg = 0
+ tvoff = 0 tvfbsdoff = 0 saref = 3E-6
+ sbref = 3E-6 wlod = 0 ku0 = -2.7E-8
+ kvsat = 0.2 kvth0 = 9.8E-9 tku0 = 0
+ llodku0 = 0 wlodku0 = 1 llodvth = 0
+ wlodvth = 1 lku0 = 0 wku0 = 0
+ pku0 = 0 lkvth0 = 0 wkvth0 = 2E-7
+ pkvth0 = 0 stk2 = 0 lodk2 = 1
+ steta0 = 0 lodeta0 = 1

.model nshort_model.19 nmos
+ level = 54 lmin = 2E-6 lmax = 4E-6 wmin = 3E-6
+ wmax = 5E-6 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 4.148E-9
+ toxm = 4.148E-9 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 9.999999999999999E22 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {2.1859E-8+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {1.1932E-8-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = 0 dwb = 0 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = 0.509180994494869 lvth0 = 4.075453062195283E-8
+ wvth0 = 4.970507576667392E-8 pvth0 = -7.846242377615352E-14 k1 = 0.539334826903307
+ lk1 = 1.75162099296683E-8 wk1 = 2.764092559425944E-9 pk1 = 1.169288997412164E-13
+ k2 = -0.024937274731741 lk2 = -1.844352958856423E-8 wk2 = -7.416269825847658E-9
+ pk2 = -1.975148544319324E-14 k3 = 2 k3b = 0.54
+ w0 = 0 lpe0 = 1.0325E-7 lpeb = -7.082E-8
+ vbm = -3 dvtp0 = 0 dvtp1 = 0
+ dvt0 = 0 dvt1 = 0.53 dvt2 = -0.032
+ dvt0w = -3.58 dvt1w = 1.6706E6 dvt2w = 0.068
+ vfbsdoff = 0 u0 = 0.03487846788479 lu0 = -8.776483274347072E-9
+ wu0 = -8.638805747076824E-9 pu0 = 1.113285114875306E-14 ua = -8.425297392492956E-10
+ lua = 2.275654349138574E-17 wua = 9.363157328877578E-16 pua = -1.640328046020571E-21
+ ub = 2.041556608872362E-18 lub = -7.780135536686935E-25 wub = -1.957190308294674E-24
+ pub = 3.392238460165525E-30 uc = 1.663509327874832E-10 luc = -1.642066561677481E-16
+ wuc = -3.226119605868081E-16 puc = 5.256731990197111E-22 ud = 0
+ up = 0 lp = 1 eu = 1.67
+ vsat = 8E4 a0 = 2.316192759607801 la0 = -3.181621248306127E-6
+ wa0 = -3.798707738142762E-6 pa0 = 1.234977999937454E-11 ags = 0.589890522317811
+ lags = -2.424929468552885E-7 wags = -1.177459808489163E-6 pags = 3.418542267468642E-12
+ b0 = 3.077719703232391E-24 lb0 = -1.223743210993162E-29 wb0 = -1.525404676617604E-29
+ pb0 = 6.065216449267613E-35 b1 = 0 keta = -0.010666299301794
+ lketa = 2.672875624490651E-8 wketa = 2.636204881437022E-8 pketa = -6.652660940626994E-14
+ a1 = 0 a2 = 0.42385546 rdsw = 65.968
+ rdswmin = 0 rdw = 0 rdwmin = 0
+ rsw = 0 rswmin = 0 prwb = 0
+ prwg = 0.021507 wr = 1 voff = -0.106555018867508
+ lvoff = 1.996499624828186E-8 wvoff = 3.057518638646371E-10 pvoff = -2.673956574776983E-14
+ voffl = 5.8197729E-9 minv = 0 nfactor = 2.291134360673405
+ lnfactor = 8.915872951937942E-7 wnfactor = 1.346086178573343E-6 pnfactor = -2.221965120692175E-12
+ eta0 = 0.274661459816246 leta0 = -7.740004381879287E-7 weta0 = -5.75474169748491E-7
+ peta0 = 2.288163563407086E-12 etab = -0.240175741331023 letab = 6.766418914329684E-7
+ wetab = 5.030874809335593E-7 petab = -2.000344244089239E-12 dsub = 1.2945715464764
+ ldsub = -2.920756370520486E-6 wdsub = -2.171600640560344E-6 pdsub = 8.634579484555043E-12
+ cit = 0 cdsc = 0 cdscb = 0
+ cdscd = 5.4E-3 pclm = 0.602364523150283 lpclm = -4.373573176073636E-7
+ wpclm = -3.800094677804715E-7 ppclm = 1.469605428271265E-12 pdiblc1 = 0.39
+ pdiblc2 = 3.244423889423422E-4 lpdiblc2 = 1.00532300833121E-8 wpdiblc2 = 5.396000589536902E-9
+ ppdiblc2 = -1.395144844266892E-14 pdiblcb = -0.025 drout = 0.56
+ pscbe1 = 7.825561224915042E8 lpscbe1 = 58.828676287745644 wpscbe1 = 75.92622305218785
+ ppscbe1 = -2.707617043800962E-4 pscbe2 = 1E-12 pvag = 0
+ delta = 0.01 fprout = 0 pdits = 0
+ pditsl = 0 pditsd = 0 lambda = 0
+ vtl = 0 lc = 5E-9 xn = 3
+ alpha0 = 3E-8 alpha1 = 0.85 beta0 = 13.86
+ aigbacc = 1 bigbacc = 0 cigbacc = 0
+ nigbacc = 0 aigbinv = 0.35 bigbinv = 0.03
+ cigbinv = 6E-3 eigbinv = 1.1 nigbinv = 0
+ aigc = 0.43 bigc = 0.054 cigc = 0.075
+ aigsd = 0.43 bigsd = 0.054 cigsd = 0.075
+ dlcig = 0 nigc = 0 poxedge = 1
+ pigcd = 1 ntox = 1 toxref = 4.148E-9
+ agidl = 0 bgidl = 2.3E9 cgidl = 0.5
+ egidl = 0.8 noia = 2.5E42 noib = 0
+ noic = 0 em = 4.1E7 af = 1
+ ef = 0.84 kf = 0 lintnoi = -1E-7
+ tnoia = 1.5E7 tnoib = 9.9E6 ntnoi = 1
+ rnoia = 0.94 rnoib = 0.26 xpart = 0
+ cgso = {2.449068E-10/sw_func_tox_lv_ratio} cgdo = {2.449068E-10/sw_func_tox_lv_ratio} cgbo = {1E-13/sw_func_tox_lv_ratio}
+ ckappas = 0.6 cf = 1.4067E-12 clc = 1E-7
+ cle = 0.6 dlc = 9.87908E-9 dwc = 0
+ vfbcv = -1 noff = 3.4037 voffcv = -0.17287
+ acde = 0.4 moin = 6.9 cgsl = {0/sw_func_tox_lv_ratio}
+ cgdl = {0/sw_func_tox_lv_ratio} ijthsrev = 0.1 ijthsfwd = 0.1
+ xjbvs = 1 bvs = 11.7 jss = 2.75E-3
+ jsws = 6E-10 cjs = {sw_nsd_pw_cj} mjs = 0.44
+ mjsws = 9E-4 cjsws = {3.67354204E-11*sw_func_nsd_pw_cj} cjswgs = {2.38232788E-10*sw_func_nsd_pw_cj}
+ mjswgs = 0.8 pbs = 0.729 pbsws = 0.2
+ pbswgs = 0.95578 xrcrg1 = 12 xrcrg2 = 1
+ rbpb = 50 rbpd = 50 rbps = 50
+ rbdb = 50 rbsb = 50 gbmin = 1E-12
+ tnom = 30 ute = -1.522233159703461 lute = -6.183638591840637E-7
+ wute = -1.229961432064954E-6 pute = 3.888438961211287E-12 kt1 = -0.295362943677519
+ lkt1 = -7.824278632453354E-8 wkt1 = -5.817825284942979E-8 pkt1 = 1.899607486602108E-13
+ kt1l = 0 kt2 = -0.040190948005096 lkt2 = -5.623986592301017E-9
+ wkt2 = -7.425247399647714E-9 pkt2 = 2.298378270937302E-14 ua1 = 1.248403605572275E-9
+ lua1 = -1.804411271650561E-15 wua1 = -3.603968215717686E-15 pua1 = 8.359019832174692E-21
+ ub1 = -1.501811367488076E-18 lub1 = 1.884257515777906E-24 wub1 = 3.569488326117102E-24
+ pub1 = -6.232784567311898E-30 uc1 = 3.168071888129177E-12 luc1 = 3.409463799904871E-17
+ wuc1 = 1.915102945280778E-17 puc1 = 1.049708130491886E-22 at = 1.619829213509008E5
+ lat = -0.087407084968485 wat = 7.745375617998557E-3 pat = -3.079666682824631E-8
+ prt = 0 njs = 1.2928 xtis = 2
+ tpb = 1.2287E-3 tpbsw = 0 tpbswg = 0
+ tcj = 7.92E-4 tcjsw = 1E-5 tcjswg = 0
+ tvoff = 0 tvfbsdoff = 0 saref = 3E-6
+ sbref = 3E-6 wlod = 0 ku0 = -2.7E-8
+ kvsat = 0.2 kvth0 = 9.8E-9 tku0 = 0
+ llodku0 = 0 wlodku0 = 1 llodvth = 0
+ wlodvth = 1 lku0 = 0 wku0 = 0
+ pku0 = 0 lkvth0 = 0 wkvth0 = 2E-7
+ pkvth0 = 0 stk2 = 0 lodk2 = 1
+ steta0 = 0 lodeta0 = 1

.model nshort_model.20 nmos
+ level = 54 lmin = 1E-6 lmax = 2E-6 wmin = 3E-6
+ wmax = 5E-6 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 4.148E-9
+ toxm = 4.148E-9 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 9.999999999999999E22 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {2.1859E-8+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {1.1932E-8-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = 0 dwb = 0 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = 0.523354715713193 lvth0 = 1.274532986845788E-8
+ wvth0 = -8.821092714134797E-8 pvth0 = 1.940783545464932E-13 k1 = 0.432298026505692
+ lk1 = 2.2903548452021E-7 wk1 = 5.852102678658033E-7 pk1 = -1.034063955344027E-12
+ k2 = 4.167122190858442E-3 lk2 = -7.595777610560314E-8 wk2 = -1.882744749270831E-7
+ pk2 = 3.376489245527416E-13 k3 = 2 k3b = 0.54
+ w0 = 0 lpe0 = 1.0325E-7 lpeb = -7.082E-8
+ vbm = -3 dvtp0 = 0 dvtp1 = 0
+ dvt0 = 0 dvt1 = 0.53 dvt2 = -0.032
+ dvt0w = -3.58 dvt1w = 1.6706E6 dvt2w = 0.068
+ vfbsdoff = 0 u0 = 0.033817816925289 lu0 = -6.680492729842284E-9
+ wu0 = -7.739682664929958E-10 pu0 = -4.409137330777942E-15 ua = -3.45811699455426E-10
+ lua = -9.588258567947126E-16 wua = 6.502986599076524E-16 pua = -1.075119411489957E-21
+ ub = 1.130976655458199E-18 lub = 1.021416273151356E-24 wub = -6.856039698890118E-25
+ pub = 8.794109197339134E-31 uc = 1.502659291625749E-10 luc = -1.324205014444364E-16
+ wuc = -2.857632556708883E-16 puc = 4.528551466819849E-22 ud = 0
+ up = 0 lp = 1 eu = 1.67
+ vsat = 6.427304154657319E4 lvsat = 0.031078608770321 wvsat = 0.059233836649858
+ pvsat = -1.17054117021903E-7 a0 = -0.610308191474134 la0 = 2.60154263516112E-6
+ wa0 = 8.041458131041097E-6 pa0 = -1.104799802069097E-11 ags = -0.421797422204469
+ lags = 1.756740021081191E-6 wags = 1.688826943756396E-6 pags = -2.245630169966887E-12
+ b0 = -6.155439406464784E-24 lb0 = 6.008546000468908E-30 wb0 = 3.050809353235209E-29
+ pb0 = -2.978004838829604E-35 b1 = 0 keta = 0.093430230494687
+ lketa = -1.789801437609941E-7 wketa = -1.258512633892627E-7 pketa = 2.342675965185683E-13
+ a1 = 0 a2 = 0.42385546 rdsw = 65.968
+ rdswmin = 0 rdw = 0 rdwmin = 0
+ rsw = 0 rswmin = 0 prwb = 0
+ prwg = 0.021507 wr = 1 voff = -0.085071212012124
+ lvoff = -2.248992789568902E-8 wvoff = 4.792095378758716E-8 pvoff = -1.208336804165071E-13
+ voffl = 5.8197729E-9 minv = 0 nfactor = 2.535915471187813
+ lnfactor = 4.078665305862956E-7 wnfactor = 2.176960982826833E-6 pnfactor = -3.86388673287045E-12
+ eta0 = -0.228774618326325 leta0 = 2.208577195284188E-7 weta0 = 1.136378996742067E-6
+ peta0 = -1.094691105608898E-12 etab = 0.081311458417059 letab = 4.133946247159329E-8
+ wetab = -4.058369249207894E-7 petab = -2.041860044018501E-13 dsub = -1.489410333773344
+ ldsub = 2.580770446388722E-6 wdsub = 6.92435486625373E-6 pdsub = -9.340265646858491E-12
+ cit = 0 cdsc = 0 cdscb = 0
+ cdscd = 5.4E-3 pclm = 1.227253434438243 lpclm = -1.672222791204307E-6
+ wpclm = -3.249432765319294E-6 ppclm = 7.139976105776442E-12 pdiblc1 = 0.22431275124467
+ lpdiblc1 = 3.274205370063626E-7 wpdiblc1 = -1.755452638519438E-7 ppdiblc1 = 3.469013155273246E-13
+ pdiblc2 = 3.212200965733015E-3 lpdiblc2 = 4.346626400407286E-9 wpdiblc2 = 9.366012296791173E-9
+ ppdiblc2 = -2.179673149779555E-14 pdiblcb = -0.049445635189418 lpdiblcb = 4.830789974067662E-8
+ wpdiblcb = 6.779777293059324E-10 ppdiblcb = -1.339776198079708E-15 drout = 0.8528408
+ ldrout = -5.786932471488001E-7 pscbe1 = 5.78453802216528E8 lpscbe1 = 462.16261906665557
+ wpscbe1 = 1.703665918007095E3 ppscbe1 = -3.487396714209506E-3 pscbe2 = 1E-12
+ pvag = 0 delta = 0.01 fprout = 0
+ pdits = 0 pditsl = 0 pditsd = 0
+ lambda = 0 vtl = 0 lc = 5E-9
+ xn = 3 alpha0 = -9.144845511177095E-6 lalpha0 = 1.813074250907545E-11
+ walpha0 = 2.70403215188267E-11 palpha0 = -5.34353528049281E-17 alpha1 = 1.086627438273912
+ lalpha1 = -4.67607999360855E-7 walpha1 = -1.337284492759069E-6 palpha1 = 2.642656028382934E-12
+ beta0 = 7.449738725241121 lbeta0 = 1.266754807445691E-5 wbeta0 = 1.701998445329724E-5
+ pbeta0 = -3.363380399760098E-11 aigbacc = 1 bigbacc = 0
+ cigbacc = 0 nigbacc = 0 aigbinv = 0.35
+ bigbinv = 0.03 cigbinv = 6E-3 eigbinv = 1.1
+ nigbinv = 0 aigc = 0.43 bigc = 0.054
+ cigc = 0.075 aigsd = 0.43 bigsd = 0.054
+ cigsd = 0.075 dlcig = 0 nigc = 0
+ poxedge = 1 pigcd = 1 ntox = 1
+ toxref = 4.148E-9 agidl = 0 bgidl = 2.3E9
+ cgidl = 0.5 egidl = 0.8 noia = 2.5E42
+ noib = 0 noic = 0 em = 4.1E7
+ af = 1 ef = 0.84 kf = 0
+ lintnoi = -1E-7 tnoia = 1.5E7 tnoib = 9.9E6
+ ntnoi = 1 rnoia = 0.94 rnoib = 0.26
+ xpart = 0 cgso = {2.449068E-10/sw_func_tox_lv_ratio} cgdo = {2.449068E-10/sw_func_tox_lv_ratio}
+ cgbo = {1E-13/sw_func_tox_lv_ratio} ckappas = 0.6 cf = 1.4067E-12
+ clc = 1E-7 cle = 0.6 dlc = 9.87908E-9
+ dwc = 0 vfbcv = -1 noff = 3.4037
+ voffcv = -0.17287 acde = 0.4 moin = 6.9
+ cgsl = {0/sw_func_tox_lv_ratio} cgdl = {0/sw_func_tox_lv_ratio} ijthsrev = 0.1
+ ijthsfwd = 0.1 xjbvs = 1 bvs = 11.7
+ jss = 2.75E-3 jsws = 6E-10 cjs = {sw_nsd_pw_cj}
+ mjs = 0.44 mjsws = 9E-4 cjsws = {3.67354204E-11*sw_func_nsd_pw_cj}
+ cjswgs = {2.38232788E-10*sw_func_nsd_pw_cj} mjswgs = 0.8 pbs = 0.729
+ pbsws = 0.2 pbswgs = 0.95578 xrcrg1 = 12
+ xrcrg2 = 1 rbpb = 50 rbpd = 50
+ rbps = 50 rbdb = 50 rbsb = 50
+ gbmin = 1E-12 tnom = 30 ute = -3.275796075280338
+ lute = 2.846914946552362E-6 wute = 3.807485546516249E-6 pute = -6.066241361254255E-12
+ kt1 = -0.367980184670481 lkt1 = 6.525875782233386E-8 wkt1 = -5.825906638624544E-8
+ pkt1 = 1.901204471995995E-13 kt1l = 0 kt2 = -0.0728232365782
+ lkt2 = 5.886185361939882E-8 wkt2 = 7.557408473254903E-8 pkt2 = -1.410341854930177E-13
+ ua1 = -2.531529433449123E-9 lua1 = 5.665250484349027E-15 wua1 = 5.963864993226372E-15
+ pua1 = -1.054831981401518E-20 ub1 = 5.4439226378042E-19 lub1 = -2.159319143302494E-24
+ wub1 = 1.901090270908001E-25 pub1 = 4.453285231487411E-31 uc1 = -1.039974793582485E-10
+ luc1 = 2.458683417768605E-16 wuc1 = 6.134067939826529E-16 puc1 = -1.069359396445761E-21
+ at = 1.771510202635417E5 lat = -0.117381311281316 wat = -0.04068308861091
+ pat = 6.490456475921246E-8 prt = 0 njs = 1.2928
+ xtis = 2 tpb = 1.2287E-3 tpbsw = 0
+ tpbswg = 0 tcj = 7.92E-4 tcjsw = 1E-5
+ tcjswg = 0 tvoff = 0 tvfbsdoff = 0
+ saref = 3E-6 sbref = 3E-6 wlod = 0
+ ku0 = -2.7E-8 kvsat = 0.2 kvth0 = 9.8E-9
+ tku0 = 0 llodku0 = 0 wlodku0 = 1
+ llodvth = 0 wlodvth = 1 lku0 = 0
+ wku0 = 0 pku0 = 0 lkvth0 = 0
+ wkvth0 = 2E-7 pkvth0 = 0 stk2 = 0
+ lodk2 = 1 steta0 = 0 lodeta0 = 1

.model nshort_model.21 nmos
+ level = 54 lmin = 5E-7 lmax = 1E-6 wmin = 3E-6
+ wmax = 5E-6 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 4.148E-9
+ toxm = 4.148E-9 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 9.999999999999999E22 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {2.1859E-8+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {1.1932E-8-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = 0 dwb = 0 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = 0.484166725129136 lvth0 = 5.09981382452175E-8
+ wvth0 = 2.621288451233161E-7 pvth0 = -1.479009093928469E-13 k1 = 0.987445294256533
+ lk1 = -3.128637488330249E-7 wk1 = -1.620513871957458E-6 pk1 = 1.119022783606493E-12
+ k2 = -0.185177382314444 lk2 = 1.08868211144185E-7 wk2 = 5.454289133267766E-7
+ pk2 = -3.785453660438279E-13 k3 = 2 k3b = 0.54
+ w0 = 0 lpe0 = 1.0325E-7 lpeb = -7.082E-8
+ vbm = -3 dvtp0 = 0 dvtp1 = 0
+ dvt0 = 0 dvt1 = 0.53 dvt2 = -0.032
+ dvt0w = -3.58 dvt1w = 1.6706E6 dvt2w = 0.068
+ vfbsdoff = 0 u0 = 0.027663267951879 lu0 = -6.728159131335937E-10
+ wu0 = -1.219950617173219E-10 pu0 = -5.04555184699485E-15 ua = -1.172891699755052E-9
+ lua = -1.514832936222369E-16 wua = -5.881447193382623E-16 pua = 1.337697549536334E-22
+ ub = 2.093119324531861E-18 lub = 8.223417673246841E-26 wub = 6.059720804876044E-25
+ pub = -3.813429597765153E-31 uc = -5.719003815159122E-11 luc = 7.008473666574451E-17
+ wuc = 3.87797601997675E-16 puc = -2.046318546791757E-22 ud = 0
+ up = 0 lp = 1 eu = 1.67
+ vsat = 7.902380490699667E4 lvsat = 0.016679857626731 wvsat = -0.153164221973937
+ pvsat = 9.027527433089376E-8 a0 = 2.58318967673665 la0 = -5.157455999226815E-7
+ wa0 = -6.396882492978076E-6 pa0 = 3.045786042676609E-12 ags = 1.407338691135728
+ lags = -2.874558805025514E-8 wags = -7.365573499132349E-7 pags = 1.218747529186111E-13
+ b0 = 0 b1 = 0 keta = -0.173803003304867
+ lketa = 8.187583614716799E-8 wketa = 3.177783144312426E-7 pketa = -1.987752050568285E-13
+ a1 = 0 a2 = 0.42385546 rdsw = 65.968
+ rdswmin = 0 rdw = 0 rdwmin = 0
+ rsw = 0 rswmin = 0 prwb = 0
+ prwg = 0.021507 wr = 1 voff = -0.077581348165335
+ lvoff = -2.980105363163857E-8 wvoff = -1.502043658417364E-7 pvoff = 7.256357658518227E-14
+ voffl = 5.8197729E-9 minv = 0 nfactor = 3.264479119037772
+ lnfactor = -3.033106743713724E-7 wnfactor = -3.97074600610832E-6 pnfactor = 2.137111376480755E-12
+ eta0 = -0.471528122612334 leta0 = 4.578181541881461E-7 weta0 = 2.91386855098321E-8
+ peta0 = -1.387397716390942E-14 etab = 0.24127872090049 letab = -1.14810341259933E-7
+ wetab = -1.198495941295101E-6 petab = 5.695569972057054E-13 dsub = 1.876654397185842
+ ldsub = -7.049665158308553E-7 wdsub = -4.975986759696901E-6 pdsub = 2.276086226530454E-12
+ cit = 0 cdsc = 0 cdscb = 0
+ cdscd = 5.4E-3 pclm = -1.38575182596622 lpclm = 8.784257116658628E-7
+ wpclm = 8.102702856269318E-6 ppclm = -3.941252151338578E-12 pdiblc1 = -0.276552881066349
+ lpdiblc1 = 8.163335118679116E-7 wpdiblc1 = 2.991574971300844E-6 ppdiblc1 = -2.744638762333777E-12
+ pdiblc2 = 9.419806540666717E-3 lpdiblc2 = -1.712840875086196E-9 wpdiblc2 = -1.199593703453638E-8
+ ppdiblc2 = -9.445637253107935E-16 pdiblcb = 0.023891270378837 lpdiblcb = -2.327889391309788E-8
+ wpdiblcb = -1.355955458611859E-9 ppdiblcb = 6.456192082416162E-16 drout = -0.249455253271172
+ ldrout = 4.972976131071086E-7 wdrout = -5.771431887499531E-7 pdrout = 5.633702436936243E-13
+ pscbe1 = 1.291806799494177E9 lpscbe1 = -234.16692228395937 wpscbe1 = -3.648774159339465E3
+ ppscbe1 = 1.737312733131255E-3 pscbe2 = 1E-12 pvag = 0
+ delta = 0.01 fprout = 0 pdits = 0
+ pditsl = 0 pditsd = 0 lambda = 0
+ vtl = 0 lc = 5E-9 xn = 3
+ alpha0 = 2.289806226154408E-5 lalpha0 = -1.314749331255751E-11 walpha0 = -7.647496507976804E-11
+ palpha0 = 4.760964499427778E-17 alpha1 = 0.376745123452176 lalpha1 = 2.253336838999744E-7
+ walpha1 = 2.674568985518137E-6 palpha1 = -1.273458578488663E-12 beta0 = 32.533291276169365
+ lbeta0 = -1.181741057839598E-5 wbeta0 = -6.304794119666078E-5 pbeta0 = 4.452338067464643E-11
+ aigbacc = 1 bigbacc = 0 cigbacc = 0
+ nigbacc = 0 aigbinv = 0.35 bigbinv = 0.03
+ cigbinv = 6E-3 eigbinv = 1.1 nigbinv = 0
+ aigc = 0.43 bigc = 0.054 cigc = 0.075
+ aigsd = 0.43 bigsd = 0.054 cigsd = 0.075
+ dlcig = 0 nigc = 0 poxedge = 1
+ pigcd = 1 ntox = 1 toxref = 4.148E-9
+ agidl = 0 bgidl = 2.3E9 cgidl = 0.5
+ egidl = 0.8 noia = 2.5E42 noib = 0
+ noic = 0 em = 4.1E7 af = 1
+ ef = 0.84 kf = 0 lintnoi = -1E-7
+ tnoia = 1.5E7 tnoib = 9.9E6 ntnoi = 1
+ rnoia = 0.94 rnoib = 0.26 xpart = 0
+ cgso = {2.449068E-10/sw_func_tox_lv_ratio} cgdo = {2.449068E-10/sw_func_tox_lv_ratio} cgbo = {1E-13/sw_func_tox_lv_ratio}
+ ckappas = 0.6 cf = 1.4067E-12 clc = 1E-7
+ cle = 0.6 dlc = 9.87908E-9 dwc = 0
+ vfbcv = -1 noff = 3.4037 voffcv = -0.17287
+ acde = 0.4 moin = 6.9 cgsl = {0/sw_func_tox_lv_ratio}
+ cgdl = {0/sw_func_tox_lv_ratio} ijthsrev = 0.1 ijthsfwd = 0.1
+ xjbvs = 1 bvs = 11.7 jss = 2.75E-3
+ jsws = 6E-10 cjs = {sw_nsd_pw_cj} mjs = 0.44
+ mjsws = 9E-4 cjsws = {3.67354204E-11*sw_func_nsd_pw_cj} cjswgs = {2.38232788E-10*sw_func_nsd_pw_cj}
+ mjswgs = 0.8 pbs = 0.729 pbsws = 0.2
+ pbswgs = 0.95578 xrcrg1 = 12 xrcrg2 = 1
+ rbpb = 50 rbpd = 50 rbps = 50
+ rbdb = 50 rbsb = 50 gbmin = 1E-12
+ tnom = 30 ute = 1.007947713174185 lute = -1.334601580134483E-6
+ wute = -6.225017667048772E-6 pute = 3.726846195622251E-12 kt1 = -0.323610722303311
+ lkt1 = 2.194812830509401E-8 wkt1 = 2.712027395281218E-7 pkt1 = -1.314790821784274E-13
+ kt1l = 0 kt2 = 9.325787445708538E-3 lkt2 = -2.13267660952031E-8
+ wkt2 = -1.304250988236091E-7 pkt2 = 6.004903354675623E-14 ua1 = 5.416821995038781E-9
+ lua1 = -2.093421485649442E-15 wua1 = -9.514190674810975E-15 pua1 = 4.560367533560124E-21
+ ub1 = -1.388221491196446E-18 lub1 = -2.728252829743963E-25 wub1 = -2.629157461873699E-24
+ pub1 = 3.197316036620591E-30 uc1 = 3.920554572110796E-10 luc1 = -2.383467875141773E-16
+ wuc1 = -1.393195215080739E-15 puc1 = 8.893570622733416E-22 at = 4.960931399346734E4
+ lat = 7.116739710329363E-3 wat = 0.100952881744091 pat = -7.335140479923683E-8
+ prt = 0 njs = 1.2928 xtis = 2
+ tpb = 1.2287E-3 tpbsw = 0 tpbswg = 0
+ tcj = 7.92E-4 tcjsw = 1E-5 tcjswg = 0
+ tvoff = 0 tvfbsdoff = 0 saref = 2.75E-6
+ sbref = 2.74E-6 wlod = 0 ku0 = -2.7E-8
+ kvsat = 0.2 kvth0 = 9.8E-9 tku0 = 0
+ llodku0 = 0 wlodku0 = 1 llodvth = 0
+ wlodvth = 1 lku0 = 0 wku0 = 0
+ pku0 = 0 lkvth0 = 0 wkvth0 = 2E-7
+ pkvth0 = 0 stk2 = 0 lodk2 = 1
+ steta0 = 0 lodeta0 = 1

.model nshort_model.22 nmos
+ level = 54 lmin = 2.5E-7 lmax = 5E-7 wmin = 3E-6
+ wmax = 5E-6 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 4.148E-9
+ toxm = 4.148E-9 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 9.999999999999999E22 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {2.1859E-8+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {1.1932E-8-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = 0 dwb = 0 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = 0.64624322953999 lvth0 = -2.617232025894919E-8
+ wvth0 = -9.127629017056416E-8 pvth0 = 2.036799810544001E-14 k1 = -0.044625814061805
+ lk1 = 1.785424603972352E-7 wk1 = 1.298853682763213E-6 pk1 = -2.709932064279886E-13
+ k2 = 0.157539365270483 lk2 = -5.431157018391182E-8 wk2 = -4.530767430230906E-7
+ pk2 = 9.687912314797237E-14 k3 = 2 k3b = 0.54
+ w0 = 0 lpe0 = 1.0325E-7 lpeb = -7.082E-8
+ vbm = -3 dvtp0 = 0 dvtp1 = 0
+ dvt0 = 0 dvt1 = 0.53 dvt2 = -0.032
+ dvt0w = -3.58 dvt1w = 1.6706E6 dvt2w = 0.068
+ vfbsdoff = 0 u0 = 0.033571049541909 lu0 = -3.485723408284328E-9
+ wu0 = -1.613181329814471E-8 pu0 = 2.577298968824742E-15 ua = -8.915624398821577E-10
+ lua = -2.854342821010772E-16 wua = -7.50981466299779E-16 pua = 2.11302192304902E-22
+ ub = 1.924065949457762E-18 lub = 1.627265745267491E-25 wub = 1.618320143145017E-25
+ pub = -1.698718852291188E-31 uc = 1.640827545044646E-10 luc = -3.527120573833927E-17
+ wuc = -2.572489332484142E-16 puc = 1.024980224267562E-22 ud = 0
+ up = 0 lp = 1 eu = 1.67
+ vsat = 1.165365893506507E5 lvsat = -1.181329507132966E-3 wvsat = -0.035306476152274
+ pvsat = 3.415895866635021E-8 a0 = 1.5 ags = 2.54768889870849
+ lags = -5.717073744831196E-7 wags = -9.153052130674594E-7 pags = 2.069830454894109E-13
+ b0 = 0 b1 = 0 keta = 0.015604950702318
+ lketa = -8.30810944199725E-9 wketa = -1.396456154669616E-7 pketa = 1.902079522918284E-14
+ a1 = 0 a2 = 0.42385546 rdsw = 65.968
+ rdswmin = 0 rdw = 0 rdwmin = 0
+ rsw = 0 rswmin = 0 prwb = 0
+ prwg = 0.021507 wr = 1 voff = -0.14001377075354
+ lvoff = -7.47296701809081E-11 wvoff = 1.676737798575887E-8 pvoff = -6.937681633866028E-15
+ voffl = 5.8197729E-9 minv = 0 nfactor = 2.495136390667723
+ lnfactor = 6.300109494382939E-8 wnfactor = 3.109409936988968E-7 pnfactor = 9.844605514054602E-14
+ eta0 = 0.49 etab = 1.910278902584502E-3 letab = -8.384087608184743E-10
+ wetab = -7.494999384690316E-9 petab = 2.47857272824996E-15 dsub = 0.315373459024082
+ ldsub = 3.841554494173266E-8 wdsub = -6.085653179816074E-7 pdsub = 1.965996509579013E-13
+ cit = 0 cdsc = 0 cdscb = 0
+ cdscd = 5.4E-3 pclm = 0.35060562644632 lpclm = 5.168341970396596E-8
+ wpclm = 3.563941331672668E-7 ppclm = -2.529557011556608E-13 pdiblc1 = 1.826620146630672
+ lpdiblc1 = -1.850628808476371E-7 wpdiblc1 = -3.000380504644126E-6 ppdiblc1 = 1.08346950160757E-13
+ pdiblc2 = 8.864730887602909E-3 lpdiblc2 = -1.448549373939008E-9 wpdiblc2 = -2.695224927837527E-8
+ ppdiblc2 = 6.176674961221678E-15 pdiblcb = -0.2924087145408 lpdiblcb = 1.273229157065983E-7
+ wpdiblcb = 1.325352998521705E-6 ppdiblcb = -6.310482753041305E-13 drout = 0.609547946542344
+ ldrout = 8.829526556070053E-8 wdrout = 1.154286377499906E-6 pdrout = -2.610257042623189E-13
+ pscbe1 = 8E8 pscbe2 = 1E-12 pvag = 0
+ delta = 0.01 fprout = 0 pdits = 0
+ pditsl = 0 pditsd = 0 lambda = 0
+ vtl = 0 lc = 5E-9 xn = 3
+ alpha0 = -1.465450644562464E-5 lalpha0 = 4.732636541398974E-12 walpha0 = 5.274076207535961E-11
+ palpha0 = -1.391461447045608E-17 alpha1 = 0.85 beta0 = -3.230690458942242
+ lbeta0 = 5.211108629033115E-6 wbeta0 = 5.985155848308522E-5 pbeta0 = -1.39934955048691E-11
+ aigbacc = 1 bigbacc = 0 cigbacc = 0
+ nigbacc = 0 aigbinv = 0.35 bigbinv = 0.03
+ cigbinv = 6E-3 eigbinv = 1.1 nigbinv = 0
+ aigc = 0.43 bigc = 0.054 cigc = 0.075
+ aigsd = 0.43 bigsd = 0.054 cigsd = 0.075
+ dlcig = 0 nigc = 0 poxedge = 1
+ pigcd = 1 ntox = 1 toxref = 4.148E-9
+ agidl = 0 bgidl = 2.3E9 cgidl = 0.5
+ egidl = 0.8 noia = 2.5E42 noib = 0
+ noic = 0 em = 4.1E7 af = 1
+ ef = 0.84 kf = 0 lintnoi = -1E-7
+ tnoia = 1.5E7 tnoib = 9.9E6 ntnoi = 1
+ rnoia = 0.94 rnoib = 0.26 xpart = 0
+ cgso = {2.449068E-10/sw_func_tox_lv_ratio} cgdo = {2.449068E-10/sw_func_tox_lv_ratio} cgbo = {1E-13/sw_func_tox_lv_ratio}
+ ckappas = 0.6 cf = 1.4067E-12 clc = 1E-7
+ cle = 0.6 dlc = 9.87908E-9 dwc = 0
+ vfbcv = -1 noff = 3.4037 voffcv = -0.17287
+ acde = 0.4 moin = 6.9 cgsl = {0/sw_func_tox_lv_ratio}
+ cgdl = {0/sw_func_tox_lv_ratio} ijthsrev = 0.1 ijthsfwd = 0.1
+ xjbvs = 1 bvs = 11.7 jss = 2.75E-3
+ jsws = 6E-10 cjs = {sw_nsd_pw_cj} mjs = 0.44
+ mjsws = 9E-4 cjsws = {3.67354204E-11*sw_func_nsd_pw_cj} cjswgs = {2.38232788E-10*sw_func_nsd_pw_cj}
+ mjswgs = 0.8 pbs = 0.729 pbsws = 0.2
+ pbswgs = 0.95578 xrcrg1 = 12 xrcrg2 = 1
+ rbpb = 50 rbpd = 50 rbps = 50
+ rbdb = 50 rbsb = 50 gbmin = 1E-12
+ tnom = 30 ute = -2.354879333079661 lute = 2.665614383606388E-7
+ wute = 6.567354299951033E-7 pute = 4.501958030081682E-13 kt1 = -0.244666596782263
+ lkt1 = -1.564001184399582E-8 wkt1 = -1.899183509902113E-7 pkt1 = 8.807726937660969E-14
+ kt1l = 0 kt2 = -0.031164523937658 lkt2 = -2.047871194372516E-9
+ wkt2 = -7.000030631214457E-8 pkt2 = 3.127861453951757E-14 ua1 = 1.356030168567833E-9
+ lua1 = -1.599323085608708E-16 wua1 = -4.530399546477231E-15 pua1 = 2.187405160879809E-21
+ ub1 = -3.727401675345551E-18 lub1 = 8.40942613185622E-25 wub1 = 1.162068865966993E-23
+ pub1 = -3.587548696306705E-30 uc1 = -3.170077007878001E-10 luc1 = 9.926370828277728E-17
+ wuc1 = 1.094375104862143E-15 puc1 = -2.95064719582982E-22 at = 9.2352465394266E4
+ lat = -0.013234813425041 wat = -0.071362710095284 pat = 8.69425183679576E-9
+ prt = 0 njs = 1.2928 xtis = 2
+ tpb = 1.2287E-3 tpbsw = 0 tpbswg = 0
+ tcj = 7.92E-4 tcjsw = 1E-5 tcjswg = 0
+ tvoff = 0 tvfbsdoff = 0 saref = 1.75E-6
+ sbref = 1.74E-6 wlod = 0 ku0 = -2.7E-8
+ kvsat = 0.2 kvth0 = 9.8E-9 tku0 = 0
+ llodku0 = 0 wlodku0 = 1 llodvth = 0
+ wlodvth = 1 lku0 = 0 wku0 = 0
+ pku0 = 0 lkvth0 = 0 wkvth0 = 2E-7
+ pkvth0 = 0 stk2 = 0 lodk2 = 1
+ steta0 = 0 lodeta0 = 1

.model nshort_model.23 nmos
+ level = 54 lmin = 1.8E-7 lmax = 2.5E-7 wmin = 3E-6
+ wmax = 5E-6 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 4.148E-9
+ toxm = 4.148E-9 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 9.999999999999999E22 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {2.1859E-8+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {1.1932E-8-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = 0 dwb = 0 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = 0.783231053860297 lvth0 = -5.715019889944595E-8
+ wvth0 = -4.870291160835884E-7 pvth0 = 1.098619591461076E-13 k1 = 0.49310500821729
+ lk1 = 5.694216317032987E-8 wk1 = -2.708135375945491E-10 pk1 = 2.27856106674908E-14
+ k2 = -0.031189443942315 lk2 = -1.163319218376653E-8 wk2 = 8.49923470717168E-8
+ pk2 = -2.479766860970697E-14 k3 = 2 k3b = 0.54
+ w0 = 0 lpe0 = 1.0325E-7 lpeb = -7.082E-8
+ vbm = -3 dvtp0 = 0 dvtp1 = 0
+ dvt0 = 0 dvt1 = 0.53 dvt2 = -0.032
+ dvt0w = -3.58 dvt1w = 1.6706E6 dvt2w = 0.068
+ vfbsdoff = 0 u0 = -4.339233702000025E-3 lu0 = 5.087156403360369E-9
+ wu0 = -1.52497420008787E-8 pu0 = 2.377830893946196E-15 ua = -6.749666626615038E-9
+ lua = 1.039293966269949E-15 wua = 7.792177347540135E-15 pua = -1.7206135692216E-21
+ ub = 7.661363530875458E-18 lub = -1.134682951344723E-24 wub = -1.347426977049325E-23
+ pub = 2.913741627980166E-30 uc = -2.264736400776449E-10 luc = 5.304765510688064E-17
+ wuc = 9.86256992764633E-16 puc = -1.787034336581303E-22 ud = 0
+ up = 0 lp = 1 eu = 1.67
+ vsat = 1.109476090866033E5 lvsat = 8.25401338576716E-5 wvsat = 0.108466938060957
+ pvsat = 1.64661386982705E-9 a0 = 1.5 ags = -2.725045681211096
+ lags = 6.206477324815758E-7 pags = 9.238183740062137E-19 b0 = 0
+ b1 = 0 keta = 7.781446191362136E-3 lketa = -6.538933425907679E-9
+ wketa = -6.967213642603057E-8 pketa = 3.197272572782876E-15 a1 = 0
+ a2 = 0.42385546 rdsw = 65.968 rdswmin = 0
+ rdw = 0 rdwmin = 0 rsw = 0
+ rswmin = 0 prwb = 0 prwg = 0.021507
+ wr = 1 voff = -0.244674014581238 lvoff = 2.359271922803934E-8
+ wvoff = 5.384288673939917E-7 pvoff = -1.249041242026861E-13 voffl = 5.8197729E-9
+ minv = 0 nfactor = -1.54058639883401 lnfactor = 9.756233036705928E-7
+ wnfactor = 1.747296422702234E-5 pnfactor = -3.782505230750284E-12 eta0 = 1.377471866503572
+ leta0 = -2.006893380036518E-7 weta0 = 6.028800405608761E-7 peta0 = -1.363328808522743E-13
+ etab = -0.035213031309549 letab = 7.556508117312647E-9 wetab = 4.354878357250671E-7
+ petab = -9.769579367213014E-14 dsub = 0.894977973601966 ldsub = -9.265390156685176E-8
+ wdsub = -1.93136380632845E-7 pdsub = 1.026562127816015E-13 cit = 0
+ cdsc = 0 cdscb = 0 cdscd = 5.225705383200001E-3
+ lcdscd = 3.941428746468453E-11 wcdscd = 1.634093419898274E-8 pcdscd = -3.69527349602116E-15
+ pclm = 0.538820676834833 lpclm = 9.121221069309148E-9 wpclm = -2.077578436770348E-7
+ ppclm = -1.253806297199978E-13 pdiblc1 = 2.35904269260067 lpdiblc1 = -3.054627857031085E-7
+ wpdiblc1 = -7.843734466953255E-6 ppdiblc1 = 1.203603641781494E-12 pdiblc2 = -0.015706087698174
+ lpdiblc2 = 4.10779725777431E-9 wpdiblc2 = 1.565499551892828E-8 ppdiblc2 = -3.458356948261357E-15
+ pdiblcb = 1.120676856473143 lpdiblcb = -1.922266029802107E-7 wpdiblcb = -4.780721519080915E-6
+ ppdiblcb = 7.497549918084555E-13 drout = 0.4516027116344 ldrout = 1.240123692018433E-7
+ wdrout = 4.896295555953786E-6 pdrout = -1.107228691841165E-12 pscbe1 = 7.850767285570925E8
+ lpscbe1 = 3.374688911013327 wpscbe1 = 100.69496085557749 ppscbe1 = -2.277075566803687E-5
+ pscbe2 = 1E-12 pvag = 0 delta = 0.01
+ fprout = 0 pdits = 0 pditsl = 0
+ pditsd = 0 lambda = 0 vtl = 0
+ lc = 5E-9 xn = 3 alpha0 = 1.083252961332164E-5
+ lalpha0 = -1.030899844826904E-12 walpha0 = -7.058061164577331E-13 palpha0 = -1.828421325831271E-18
+ alpha1 = 1.837382487856127 lalpha1 = -2.23282726273833E-7 walpha1 = -2.918981075964286E-6
+ palpha1 = 6.600867045942596E-13 beta0 = 9.327764020210857 lbeta0 = 2.371189966935348E-6
+ wbeta0 = 6.112838551307019E-5 pbeta0 = -1.428223206212178E-11 aigbacc = 1
+ bigbacc = 0 cigbacc = 0 nigbacc = 0
+ aigbinv = 0.35 bigbinv = 0.03 cigbinv = 6E-3
+ eigbinv = 1.1 nigbinv = 0 aigc = 0.43
+ bigc = 0.054 cigc = 0.075 aigsd = 0.43
+ bigsd = 0.054 cigsd = 0.075 dlcig = 0
+ nigc = 0 poxedge = 1 pigcd = 1
+ ntox = 1 toxref = 4.148E-9 agidl = 0
+ bgidl = 2.3E9 cgidl = 0.5 egidl = 0.8
+ noia = 2.5E42 noib = 0 noic = 0
+ em = 4.1E7 af = 1 ef = 0.84
+ kf = 0 lintnoi = -1E-7 tnoia = 1.5E7
+ tnoib = 9.9E6 ntnoi = 1 rnoia = 0.94
+ rnoib = 0.26 xpart = 0 cgso = {2.449068E-10/sw_func_tox_lv_ratio}
+ cgdo = {2.449068E-10/sw_func_tox_lv_ratio} cgbo = {1E-13/sw_func_tox_lv_ratio} ckappas = 0.6
+ cf = 1.4067E-12 clc = 1E-7 cle = 0.6
+ dlc = 9.87908E-9 dwc = 0 vfbcv = -1
+ noff = 3.4037 voffcv = -0.17287 acde = 0.4
+ moin = 6.9 cgsl = {0/sw_func_tox_lv_ratio} cgdl = {0/sw_func_tox_lv_ratio}
+ ijthsrev = 0.1 ijthsfwd = 0.1 xjbvs = 1
+ bvs = 11.7 jss = 2.75E-3 jsws = 6E-10
+ cjs = {sw_nsd_pw_cj} mjs = 0.44 mjsws = 9E-4
+ cjsws = {3.67354204E-11*sw_func_nsd_pw_cj} cjswgs = {2.38232788E-10*sw_func_nsd_pw_cj} mjswgs = 0.8
+ pbs = 0.729 pbsws = 0.2 pbswgs = 0.95578
+ xrcrg1 = 12 xrcrg2 = 1 rbpb = 50
+ rbpd = 50 rbps = 50 rbdb = 50
+ rbsb = 50 gbmin = 1E-12 tnom = 30
+ ute = 1.987849025771341 lute = -7.154857817964913E-7 wute = 1.418809837385944E-7
+ pute = 5.666229280668301E-13 kt1 = -0.333190606036723 lkt1 = 4.378453512770768E-9
+ wkt1 = 2.874000946892423E-7 pkt1 = -1.986161465555926E-14 kt1l = 0
+ kt2 = -0.026506558540585 lkt2 = -3.101204857405105E-9 wkt2 = 1.053719628605378E-7
+ pkt2 = -8.379368922116127E-15 ua1 = 5.008738400211296E-9 lua1 = -9.859411372317968E-16
+ wua1 = 8.159284493457703E-15 pua1 = -6.821892291749174E-22 ub1 = -2.016597456236565E-18
+ lub1 = 4.540681902931925E-25 wub1 = -1.249786235522677E-23 pub1 = 1.866523955997973E-30
+ uc1 = 3.321514217833871E-10 luc1 = -4.753453905898066E-17 wuc1 = -1.467657293894471E-15
+ puc1 = 2.843030389422436E-22 at = 1.150888746399687E5 lat = -0.018376334066228
+ wat = -0.622818723869302 pat = 1.33398308967597E-7 prt = 0
+ njs = 1.2928 xtis = 2 tpb = 1.2287E-3
+ tpbsw = 0 tpbswg = 0 tcj = 7.92E-4
+ tcjsw = 1E-5 tcjswg = 0 tvoff = 0
+ tvfbsdoff = 0 saref = 1.25E-6 sbref = 1.24E-6
+ wlod = 0 ku0 = -2.7E-8 kvsat = 0.2
+ kvth0 = 9.8E-9 tku0 = 0 llodku0 = 0
+ wlodku0 = 1 llodvth = 0 wlodvth = 1
+ lku0 = 0 wku0 = 0 pku0 = 0
+ lkvth0 = 0 wkvth0 = 2E-7 pkvth0 = 0
+ stk2 = 0 lodk2 = 1 steta0 = 0
+ lodeta0 = 1

.model nshort_model.24 nmos
+ level = 54 lmin = 1.5E-7 lmax = 1.8E-7 wmin = 3E-6
+ wmax = 5E-6 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 4.148E-9
+ toxm = 4.148E-9 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 9.999999999999999E22 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {2.1859E-8+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {1.1932E-8-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = 0 dwb = 0 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = 0.530486024164743 lvth0 = -1.768760094290095E-8
+ wvth0 = 5.131328280677948E-7 pvth0 = -4.629932616591278E-14 k1 = 0.706907426128423
+ lk1 = 2.355990884735716E-8 wk1 = 5.917473316343934E-7 pk1 = -6.96497344470827E-14
+ k2 = -0.100511325281607 lk2 = -8.095509189748102E-10 wk2 = -9.690911798949731E-8
+ pk2 = 3.603698539090753E-15 k3 = 2 k3b = 0.54
+ w0 = 0 lpe0 = 1.0325E-7 lpeb = -7.082E-8
+ vbm = -3 dvtp0 = 0 dvtp1 = 0
+ dvt0 = 0 dvt1 = 0.53 dvt2 = -0.032
+ dvt0w = -3.58 dvt1w = 1.6706E6 dvt2w = 0.068
+ vfbsdoff = 0 u0 = 0.163526774867455 lu0 = -2.112277071064005E-8
+ wu0 = -3.762372092908162E-7 pu0 = 5.874097008672789E-14 ua = 1.697280683153368E-8
+ lua = -2.664638149591559E-15 wua = -5.375949692198014E-14 pua = 7.889818644524217E-21
+ ub = -1.396242758100361E-17 lub = 2.241569297699627E-24 wub = 5.054657819396402E-23
+ pub = -7.082217489798333E-30 uc = 5.266491414273811E-10 luc = -6.454192350618809E-17
+ wuc = -1.380318046719221E-15 puc = 1.908041267067207E-22 ud = 0
+ up = 0 lp = 1 eu = 1.67
+ vsat = -9.405219097907498E4 lvsat = 0.032090388916912 wvsat = 0.549261948091962
+ pvsat = -6.717735581637394E-8 a0 = 1.5 ags = 1.25
+ b0 = 0 b1 = 0 keta = 0.551933959366785
+ lketa = -9.150073022306555E-8 wketa = -2.6412779467076E-6 pketa = 4.04717517366906E-13
+ a1 = 0 a2 = 0.42385546 rdsw = 65.968
+ rdswmin = 0 rdw = 0 rdwmin = 0
+ rsw = 0 rswmin = 0 prwb = 0
+ prwg = 0.021507 wr = 1 voff = 0.09710513753736
+ lvoff = -2.977131046715003E-8 wvoff = -8.252317454892215E-7 pvoff = 8.801238925044721E-14
+ voffl = 5.8197729E-9 minv = 0 nfactor = 9.877720444576628
+ lnfactor = -8.071854536321703E-7 wnfactor = -3.245888202100074E-5 pnfactor = 4.013653515031048E-12
+ eta0 = 0.476332994046942 leta0 = -5.998911901376343E-8 weta0 = -1.406122567555263E-6
+ peta0 = 1.773447503685473E-13 etab = 0.150032677917453 letab = -2.136701593855456E-8
+ wetab = -5.947852485411629E-7 petab = 6.316692461286194E-14 dsub = 0.328974217717204
+ ldsub = -4.280339138028589E-9 wdsub = 3.833604585024334E-7 pdsub = 1.264430230637563E-14
+ cit = 0 cdsc = 0 cdscb = 0
+ cdscd = 5.254590318563202E-3 lcdscd = 3.490430919681573E-11 wcdscd = 5.118232552580531E-9
+ pcdscd = -1.943005751758505E-15 pclm = 2.605040017659816 lpclm = -3.134900019297404E-7
+ wpclm = -5.75625340065393E-6 ppclm = 7.409392725641468E-13 pdiblc1 = 0.731199149596757
+ lpdiblc1 = -5.129780627264961E-8 wpdiblc1 = -1.1063205428219E-6 ppdiblc1 = 1.516507813233211E-13
+ pdiblc2 = 0.014626832942761 lpdiblc2 = -6.282636394187536E-10 wpdiblc2 = -1.839020505447893E-8
+ ppdiblc2 = 1.857324488468152E-15 pdiblcb = -0.843678184823999 lpdiblcb = 1.144799357477598E-7
+ wpdiblcb = 2.188779206060721E-6 ppdiblcb = -3.384349734122589E-13 drout = 4.635200134652515
+ ldrout = -5.291977980385129E-7 wdrout = -1.221498317939268E-5 pdrout = 1.564457924780891E-12
+ pscbe1 = 8.624336048959348E8 lpscbe1 = -8.703504333028153 wpscbe1 = -209.93659666280394
+ ppscbe1 = 2.573001319665313E-5 pscbe2 = 1E-12 pvag = 0
+ delta = 0.01 fprout = 0 pdits = 0
+ pditsl = 0 pditsd = 0 lambda = 0
+ vtl = 0 lc = 5E-9 xn = 3
+ alpha0 = 2.188879729595615E-5 lalpha0 = -2.757181255722723E-12 walpha0 = -6.462076898768381E-11
+ palpha0 = 8.151005317030483E-18 alpha1 = -1.453892471664294 lalpha1 = 2.906037808058473E-7
+ walpha1 = 6.81095584391666E-6 palpha1 = -8.591067263282717E-13 beta0 = 69.31149233316634
+ lbeta0 = -6.99442943693627E-6 wbeta0 = -1.579296820551016E-4 pbeta0 = 1.99206183757023E-11
+ aigbacc = 1 bigbacc = 0 cigbacc = 0
+ nigbacc = 0 aigbinv = 0.35 bigbinv = 0.03
+ cigbinv = 6E-3 eigbinv = 1.1 nigbinv = 0
+ aigc = 0.43 bigc = 0.054 cigc = 0.075
+ aigsd = 0.43 bigsd = 0.054 cigsd = 0.075
+ dlcig = 0 nigc = 0 poxedge = 1
+ pigcd = 1 ntox = 1 toxref = 4.148E-9
+ agidl = 0 bgidl = 2.3E9 cgidl = 0.5
+ egidl = 0.8 noia = 2.5E42 noib = 0
+ noic = 0 em = 4.1E7 af = 1
+ ef = 0.84 kf = 0 lintnoi = -1E-7
+ tnoia = 1.5E7 tnoib = 9.9E6 ntnoi = 1
+ rnoia = 0.94 rnoib = 0.26 xpart = 0
+ cgso = {2.449068E-10/sw_func_tox_lv_ratio} cgdo = {2.449068E-10/sw_func_tox_lv_ratio} cgbo = {1E-13/sw_func_tox_lv_ratio}
+ ckappas = 0.6 cf = 1.4067E-12 clc = 1E-7
+ cle = 0.6 dlc = 9.87908E-9 dwc = 0
+ vfbcv = -1 noff = 3.4037 voffcv = -0.17287
+ acde = 0.4 moin = 6.9 cgsl = {0/sw_func_tox_lv_ratio}
+ cgdl = {0/sw_func_tox_lv_ratio} ijthsrev = 0.1 ijthsfwd = 0.1
+ xjbvs = 1 bvs = 11.7 jss = 2.75E-3
+ jsws = 6E-10 cjs = {sw_nsd_pw_cj} mjs = 0.44
+ mjsws = 9E-4 cjsws = {3.67354204E-11*sw_func_nsd_pw_cj} cjswgs = {2.38232788E-10*sw_func_nsd_pw_cj}
+ mjswgs = 0.8 pbs = 0.729 pbsws = 0.2
+ pbswgs = 0.95578 xrcrg1 = 12 xrcrg2 = 1
+ rbpb = 50 rbpd = 50 rbps = 50
+ rbdb = 50 rbsb = 50 gbmin = 1E-12
+ tnom = 30 ute = -21.701412033642193 lute = 2.9832606829761E-6
+ wute = 6.02560301002574E-5 pute = -8.819359858389951E-12 kt1 = -0.642586378648221
+ lkt1 = 5.268627186523972E-8 wkt1 = 1.157755826274241E-6 pkt1 = -1.557554771623146E-13
+ kt1l = 0 kt2 = -0.116745068188598 lkt2 = 1.098827508499715E-8
+ wkt2 = 2.597570561299275E-7 pkt2 = -3.248443984482556E-14 ua1 = -2.58429561152692E-8
+ lua1 = 3.831119037637265E-15 wua1 = 7.632856654019548E-14 pua1 = -1.132586825082437E-20
+ ub1 = 1.540697490159957E-17 lub1 = -2.266378703369911E-24 wub1 = -4.345504461913664E-23
+ pub1 = 6.700054565955806E-30 uc1 = -4.011452665842779E-10 luc1 = 6.695947267599305E-17
+ wuc1 = 1.621022592510802E-15 puc1 = -1.979510838015301E-22 at = -2.489356391281495E5
+ lat = 0.038460997415471 wat = 1.146221855038378 pat = -1.428126108607324E-7
+ prt = 0 njs = 1.2928 xtis = 2
+ tpb = 1.2287E-3 tpbsw = 0 tpbswg = 0
+ tcj = 7.92E-4 tcjsw = 1E-5 tcjswg = 0
+ tvoff = 0 tvfbsdoff = 0 saref = 1.1E-6
+ sbref = 1.1E-6 wlod = 0 ku0 = -2.7E-8
+ kvsat = 0.2 kvth0 = 9.8E-9 tku0 = 0
+ llodku0 = 0 wlodku0 = 1 llodvth = 0
+ wlodvth = 1 lku0 = 0 wku0 = 0
+ pku0 = 0 lkvth0 = 0 wkvth0 = 2E-7
+ pkvth0 = 0 stk2 = 0 lodk2 = 1
+ steta0 = 0 lodeta0 = 1

.model nshort_model.25 nmos
+ level = 54 lmin = 8E-6 lmax = 2.02E-5 wmin = 1E-6
+ wmax = 3E-6 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 4.148E-9
+ toxm = 4.148E-9 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 9.999999999999999E22 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {2.1859E-8+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {1.1932E-8-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = 0 dwb = 0 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = 0.5190122089033 wvth0 = 7.744250006534551E-9
+ k1 = 0.58873918469163 wk1 = -1.101858766289213E-7 k2 = -0.044527264341045
+ wk2 = 4.337667538500889E-8 k3 = 2 k3b = 0.54
+ w0 = 0 lpe0 = 1.0325E-7 lpeb = -7.082E-8
+ vbm = -3 dvtp0 = 0 dvtp1 = 0
+ dvt0 = 0 dvt1 = 0.53 dvt2 = -0.032
+ dvt0w = -3.58 dvt1w = 1.6706E6 dvt2w = 0.068
+ vfbsdoff = 0 u0 = 0.0319277721535 wu0 = -3.199501686493289E-9
+ ua = -7.2528366620603E-10 wua = 6.062561670793479E-17 ub = 1.625898568659E-18
+ wub = -2.470818181123657E-25 uc = 9.257106339300001E-11 wuc = -6.385292232558483E-17
+ ud = 0 up = 0 lp = 1
+ eu = 1.67 vsat = 8E4 a0 = 1.450186822348
+ wa0 = -8.258912504459001E-8 ags = 0.448590173269 wags = -9.895909590002584E-8
+ b0 = 3.1148865293E-24 wb0 = -2.978709920012062E-30 b1 = 0
+ keta = -7.6300127798643E-3 wketa = 5.830121513082793E-9 a1 = 0
+ a2 = 0.42385546 rdsw = 65.968 rdswmin = 0
+ rdw = 0 rdwmin = 0 rsw = 0
+ rswmin = 0 prwb = 0 prwg = 0.021507
+ wr = 1 voff = -0.1030376408569 wvoff = -8.013384144421948E-9
+ voffl = 5.8197729E-9 minv = 0 nfactor = 2.61563341875
+ wnfactor = 2.915384240509128E-7 eta0 = 0.08 etab = -0.07
+ dsub = 0.56 cit = 0 cdsc = 0
+ cdscb = 0 cdscd = 5.4E-3 pclm = 0.083531
+ pdiblc1 = 0.39 pdiblc2 = 2.1336549940086E-3 wpdiblc2 = 9.722688413208678E-10
+ pdiblcb = -2.6517431834214 wpdiblcb = 4.142536962901834E-7 drout = 0.56
+ pscbe1 = 8.0881723871918E8 wpscbe1 = -45.23542698525488 pscbe2 = 1E-12
+ pvag = 0 delta = 0.01 fprout = 0
+ pdits = 0 pditsl = 0 pditsd = 0
+ lambda = 0 vtl = 0 lc = 5E-9
+ xn = 3 alpha0 = 3E-8 alpha1 = 0.85
+ beta0 = 13.86 aigbacc = 1 bigbacc = 0
+ cigbacc = 0 nigbacc = 0 aigbinv = 0.35
+ bigbinv = 0.03 cigbinv = 6E-3 eigbinv = 1.1
+ nigbinv = 0 aigc = 0.43 bigc = 0.054
+ cigc = 0.075 aigsd = 0.43 bigsd = 0.054
+ cigsd = 0.075 dlcig = 0 nigc = 0
+ poxedge = 1 pigcd = 1 ntox = 1
+ toxref = 4.148E-9 agidl = 0 bgidl = 2.3E9
+ cgidl = 0.5 egidl = 0.8 noia = 2.5E42
+ noib = 0 noic = 0 em = 4.1E7
+ af = 1 ef = 0.84 kf = 0
+ lintnoi = -1E-7 tnoia = 1.5E7 tnoib = 9.9E6
+ ntnoi = 1 rnoia = 0.94 rnoib = 0.26
+ xpart = 0 cgso = {2.449068E-10/sw_func_tox_lv_ratio} cgdo = {2.449068E-10/sw_func_tox_lv_ratio}
+ cgbo = {1E-13/sw_func_tox_lv_ratio} ckappas = 0.6 cf = 1.4067E-12
+ clc = 1E-7 cle = 0.6 dlc = 9.87908E-9
+ dwc = 0 vfbcv = -1 noff = 3.4037
+ voffcv = -0.17287 acde = 0.4 moin = 6.9
+ cgsl = {0/sw_func_tox_lv_ratio} cgdl = {0/sw_func_tox_lv_ratio} ijthsrev = 0.1
+ ijthsfwd = 0.1 xjbvs = 1 bvs = 11.7
+ jss = 2.75E-3 jsws = 6E-10 cjs = {sw_nsd_pw_cj}
+ mjs = 0.44 mjsws = 9E-4 cjsws = {3.67354204E-11*sw_func_nsd_pw_cj}
+ cjswgs = {2.38232788E-10*sw_func_nsd_pw_cj} mjswgs = 0.8 pbs = 0.729
+ pbsws = 0.2 pbswgs = 0.95578 xrcrg1 = 12
+ xrcrg2 = 1 rbpb = 50 rbpd = 50
+ rbps = 50 rbdb = 50 rbsb = 50
+ gbmin = 1E-12 tnom = 30 ute = -2.0306136666
+ wute = 7.10434966923581E-7 kt1 = -0.32774844426 wkt1 = 3.37265784138413E-8
+ kt1l = 0 kt2 = -0.050827695750128 wkt2 = 2.88711497868959E-8
+ ua1 = -1.581243635199999E-10 wua1 = 1.445634797795632E-15 ub1 = -1.780089171E-19
+ wub1 = -7.306482976577779E-25 uc1 = 3.4090075257355E-11 wuc1 = -5.594096528233995E-17
+ at = 1.4E5 prt = 0 njs = 1.2928
+ xtis = 2 tpb = 1.2287E-3 tpbsw = 0
+ tpbswg = 0 tcj = 7.92E-4 tcjsw = 1E-5
+ tcjswg = 0 tvoff = 0 tvfbsdoff = 0
+ saref = 3E-6 sbref = 3E-6 wlod = 0
+ ku0 = -2.7E-8 kvsat = 0.2 kvth0 = 9.8E-9
+ tku0 = 0 llodku0 = 0 wlodku0 = 1
+ llodvth = 0 wlodvth = 1 lku0 = 0
+ wku0 = 0 pku0 = 0 lkvth0 = 0
+ wkvth0 = 2E-7 pkvth0 = 0 stk2 = 0
+ lodk2 = 1 steta0 = 0 lodeta0 = 1

.model nshort_model.26 nmos
+ level = 54 lmin = 4E-6 lmax = 8E-6 wmin = 1E-6
+ wmax = 3E-6 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 4.148E-9
+ toxm = 4.148E-9 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 9.999999999999999E22 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {2.1859E-8+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {1.1932E-8-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = 0 dwb = 0 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = 0.509638935233853 lvth0 = 7.476250555272892E-8
+ wvth0 = 1.212938469420435E-8 pvth0 = -3.497643064717184E-14 k1 = 0.592058106662426
+ lk1 = -2.64721730124561E-8 wk1 = -1.292697343703535E-7 pk1 = 1.522154447503158E-13
+ k2 = -0.042850132665813 lk2 = -1.337703033155827E-8 wk2 = 4.990943417686033E-8
+ pk2 = -5.210617257900274E-14 k3 = 2 k3b = 0.54
+ w0 = 0 lpe0 = 1.0325E-7 lpeb = -7.082E-8
+ vbm = -3 dvtp0 = 0 dvtp1 = 0
+ dvt0 = 0 dvt1 = 0.53 dvt2 = -0.032
+ dvt0w = -3.58 dvt1w = 1.6706E6 dvt2w = 0.068
+ vfbsdoff = 0 u0 = 0.031831364715018 lu0 = 7.6895884074524E-10
+ wu0 = -2.47546057509716E-9 pu0 = -5.775050374086675E-15 ua = -8.093546335486154E-10
+ lua = 6.705614691760204E-16 wua = 1.765052421675274E-16 pua = -9.242716522947734E-22
+ ub = 1.732026797736255E-18 lub = -8.464931885593393E-25 wub = -3.554449048445456E-25
+ pub = 8.643187171556622E-31 uc = 1.075427148975038E-10 luc = -1.194159285445268E-16
+ wuc = -7.77688997509046E-17 puc = 1.109957285172802E-22 ud = 0
+ up = 0 lp = 1 eu = 1.67
+ vsat = 8E4 a0 = 1.595203041198602 la0 = -1.156669083758166E-6
+ wa0 = -9.823616912863295E-8 pa0 = 1.248029516123218E-13 ags = 0.435165442136222
+ lags = 1.070774812784697E-7 wags = -7.785314996873841E-8 pags = -1.68343895156595E-13
+ b0 = 6.211189645566196E-24 lb0 = -2.4696534752563E-29 wb0 = -5.939648856641333E-30
+ pb0 = 2.361685164625044E-35 b1 = 0 keta = -9.567200954886874E-3
+ lketa = 1.545127634157186E-8 wketa = -3.052653003699155E-9 pketa = 7.08502176031871E-14
+ a1 = 0 a2 = 0.42385546 rdsw = 65.968
+ rdswmin = 0 rdw = 0 rdwmin = 0
+ rsw = 0 rswmin = 0 prwb = 0
+ prwg = 0.021507 wr = 1 voff = -0.103469589465304
+ lvoff = 3.445280845639406E-9 wvoff = -1.274024993766634E-8 pvoff = 3.770212442066515E-14
+ voffl = 5.8197729E-9 minv = 0 nfactor = 2.502740809060162
+ lnfactor = 9.004468082810604E-7 wnfactor = 4.271573801385408E-7 pnfactor = -1.081715237932948E-12
+ eta0 = 0.08 etab = -0.07 dsub = 0.56
+ cit = 0 cdsc = 0 cdscb = 0
+ cdscd = 5.4E-3 pclm = -0.298309837363718 lpclm = 3.045614449166896E-6
+ wpclm = -6.225938607793996E-8 ppclm = 4.965893306341557E-13 pdiblc1 = 0.39
+ pdiblc2 = 7.145437056862555E-4 lpdiblc2 = 1.131902463479423E-8 wpdiblc2 = 2.144671813787257E-9
+ ppdiblc2 = -9.35124555519617E-15 pdiblcb = -5.262815217010509 lpdiblcb = 2.08262656457033E-5
+ wpdiblcb = 8.260359550282996E-7 ppdiblcb = -3.284431298082403E-12 drout = 0.56
+ pscbe1 = 7.915496146003578E8 lpscbe1 = 137.72891836860597 wpscbe1 = -13.242280145052295
+ ppscbe1 = -2.551816902654261E-4 pscbe2 = 1E-12 pvag = 0
+ delta = 0.01 fprout = 0 pdits = 0
+ pditsl = 0 pditsd = 0 lambda = 0
+ vtl = 0 lc = 5E-9 xn = 3
+ alpha0 = 3E-8 alpha1 = 0.85 beta0 = 13.86
+ aigbacc = 1 bigbacc = 0 cigbacc = 0
+ nigbacc = 0 aigbinv = 0.35 bigbinv = 0.03
+ cigbinv = 6E-3 eigbinv = 1.1 nigbinv = 0
+ aigc = 0.43 bigc = 0.054 cigc = 0.075
+ aigsd = 0.43 bigsd = 0.054 cigsd = 0.075
+ dlcig = 0 nigc = 0 poxedge = 1
+ pigcd = 1 ntox = 1 toxref = 4.148E-9
+ agidl = 0 bgidl = 2.3E9 cgidl = 0.5
+ egidl = 0.8 noia = 2.5E42 noib = 0
+ noic = 0 em = 4.1E7 af = 1
+ ef = 0.84 kf = 0 lintnoi = -1E-7
+ tnoia = 1.5E7 tnoib = 9.9E6 ntnoi = 1
+ rnoia = 0.94 rnoib = 0.26 xpart = 0
+ cgso = {2.449068E-10/sw_func_tox_lv_ratio} cgdo = {2.449068E-10/sw_func_tox_lv_ratio} cgbo = {1E-13/sw_func_tox_lv_ratio}
+ ckappas = 0.6 cf = 1.4067E-12 clc = 1E-7
+ cle = 0.6 dlc = 9.87908E-9 dwc = 0
+ vfbcv = -1 noff = 3.4037 voffcv = -0.17287
+ acde = 0.4 moin = 6.9 cgsl = {0/sw_func_tox_lv_ratio}
+ cgdl = {0/sw_func_tox_lv_ratio} ijthsrev = 0.1 ijthsfwd = 0.1
+ xjbvs = 1 bvs = 11.7 jss = 2.75E-3
+ jsws = 6E-10 cjs = {sw_nsd_pw_cj} mjs = 0.44
+ mjsws = 9E-4 cjsws = {3.67354204E-11*sw_func_nsd_pw_cj} cjswgs = {2.38232788E-10*sw_func_nsd_pw_cj}
+ mjswgs = 0.8 pbs = 0.729 pbsws = 0.2
+ pbswgs = 0.95578 xrcrg1 = 12 xrcrg2 = 1
+ rbpb = 50 rbpd = 50 rbps = 50
+ rbdb = 50 rbsb = 50 gbmin = 1E-12
+ tnom = 30 ute = -1.974622851752129 lute = -4.465903539774344E-7
+ wute = 4.64685325194136E-7 pute = 1.960132564385329E-12 kt1 = -0.325071153253314
+ lkt1 = -2.135443718090489E-8 wkt1 = 3.23355427059388E-8 pkt1 = 1.109508998708666E-14
+ kt1l = 0 kt2 = -0.049240629398559 lkt2 = -1.265865706113848E-8
+ wkt2 = 2.741214020582045E-8 pkt2 = 1.16372588439608E-14 ua1 = -4.468090853822071E-11
+ lua1 = -9.048404252445485E-16 wua1 = 1.240287085658929E-15 pua1 = 1.637881279291194E-21
+ ub1 = -2.903103558939177E-19 lub1 = 8.957315488159626E-25 wub1 = -6.173533711029913E-25
+ pub1 = -9.036557423109887E-31 uc1 = 1.939238192629858E-11 luc1 = 1.17230800894799E-16
+ wuc1 = -4.770669428224664E-17 puc1 = -6.567766535760025E-23 at = 1.4E5
+ prt = 0 njs = 1.2928 xtis = 2
+ tpb = 1.2287E-3 tpbsw = 0 tpbswg = 0
+ tcj = 7.92E-4 tcjsw = 1E-5 tcjswg = 0
+ tvoff = 0 tvfbsdoff = 0 saref = 3E-6
+ sbref = 3E-6 wlod = 0 ku0 = -2.7E-8
+ kvsat = 0.2 kvth0 = 9.8E-9 tku0 = 0
+ llodku0 = 0 wlodku0 = 1 llodvth = 0
+ wlodvth = 1 lku0 = 0 wku0 = 0
+ pku0 = 0 lkvth0 = 0 wkvth0 = 2E-7
+ pkvth0 = 0 stk2 = 0 lodk2 = 1
+ steta0 = 0 lodeta0 = 1

.model nshort_model.27 nmos
+ level = 54 lmin = 2E-6 lmax = 4E-6 wmin = 1E-6
+ wmax = 3E-6 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 4.148E-9
+ toxm = 4.148E-9 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 9.999999999999999E22 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {2.1859E-8+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {1.1932E-8-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = 0 dwb = 0 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = 0.533942027629884 lvth0 = -2.186989503445662E-8
+ wvth0 = -2.349552079177494E-8 pvth0 = 1.066730385522279E-13 k1 = 0.587413998701035
+ lk1 = -8.006568159283508E-9 wk1 = -1.393714976011039E-7 pk1 = 1.92381429195579E-13
+ k2 = -0.048536277524039 lk2 = 9.231854940448377E-9 wk2 = 6.234903734697046E-8
+ pk2 = -1.015677265693917E-13 k3 = 2 k3b = 0.54
+ w0 = 0 lpe0 = 1.0325E-7 lpeb = -7.082E-8
+ vbm = -3 dvtp0 = 0 dvtp1 = 0
+ dvt0 = 0 dvt1 = 0.53 dvt2 = -0.032
+ dvt0w = -3.58 dvt1w = 1.6706E6 dvt2w = 0.068
+ vfbsdoff = 0 u0 = 0.033253834963507 lu0 = -4.886976323199988E-9
+ wu0 = -3.835932685278684E-9 pu0 = -3.656282397979482E-16 ua = -6.58944617912882E-10
+ lua = 7.251079124621755E-17 wua = 3.93586343213102E-16 pua = -1.78741563308172E-21
+ ub = 1.645880168214199E-18 lub = -5.039624736380313E-25 wub = -7.87459168952881E-25
+ pub = 2.582066185190323E-30 uc = 8.601730917956173E-11 luc = -3.382798795481161E-17
+ wuc = -8.512311511993483E-17 puc = 1.402370889978347E-22 ud = 0
+ up = 0 lp = 1 eu = 1.67
+ vsat = 8E4 a0 = 0.841633167379816 la0 = 1.839627220048167E-6
+ wa0 = 5.605062422881676E-7 pa0 = -2.49444646514883E-12 ags = 0.198529086458479
+ lags = 1.047975813997548E-6 wags = -2.048504016406662E-8 pags = -3.964473018029036E-13
+ b0 = -3.07771970323239E-24 lb0 = 1.223743210993163E-29 wb0 = 2.943167953246477E-30
+ pb0 = -1.170243605294964E-35 b1 = 0 keta = -0.016040764210479
+ lketa = 4.119104425040748E-8 wketa = 4.225048268354481E-8 pketa = -1.092812111157484E-13
+ a1 = 0 a2 = 0.42385546 rdsw = 65.968
+ rdswmin = 0 rdw = 0 rdwmin = 0
+ rsw = 0 rswmin = 0 prwb = 0
+ prwg = 0.021507 wr = 1 voff = -0.116034829726726
+ lvoff = 5.340638499772913E-8 wvoff = 2.833074607037478E-8 pvoff = -1.256017413627634E-13
+ voffl = 5.8197729E-9 minv = 0 nfactor = 2.441503227177515
+ lnfactor = 1.143935762157604E-6 wnfactor = 9.015534051668424E-7 pnfactor = -2.96797835130488E-12
+ eta0 = 0.08 etab = -0.07 dsub = 0.56
+ cit = 0 cdsc = 0 cdscb = 0
+ cdscd = 5.4E-3 pclm = 0.456754698374247 lpclm = 4.33751662958847E-8
+ wpclm = 5.045423622807617E-8 ppclm = 4.842463929280194E-14 pdiblc1 = 0.39
+ pdiblc2 = 2.500686019538757E-3 lpdiblc2 = 4.217079879561998E-9 wpdiblc2 = -1.03758928320993E-9
+ ppdiblc2 = 3.301857353973834E-15 pdiblcb = -0.025 drout = 0.56
+ pscbe1 = 8.642431193654155E8 lpscbe1 = -151.31034289391135 wpscbe1 = -165.5635754402125
+ ppscbe1 = 3.50468495524291E-4 pscbe2 = 1E-12 pvag = 0
+ delta = 0.01 fprout = 0 pdits = 0
+ pditsl = 0 pditsd = 0 lambda = 0
+ vtl = 0 lc = 5E-9 xn = 3
+ alpha0 = 3E-8 alpha1 = 0.85 beta0 = 13.86
+ aigbacc = 1 bigbacc = 0 cigbacc = 0
+ nigbacc = 0 aigbinv = 0.35 bigbinv = 0.03
+ cigbinv = 6E-3 eigbinv = 1.1 nigbinv = 0
+ aigc = 0.43 bigc = 0.054 cigc = 0.075
+ aigsd = 0.43 bigsd = 0.054 cigsd = 0.075
+ dlcig = 0 nigc = 0 poxedge = 1
+ pigcd = 1 ntox = 1 toxref = 4.148E-9
+ agidl = 0 bgidl = 2.3E9 cgidl = 0.5
+ egidl = 0.8 noia = 2.5E42 noib = 0
+ noic = 0 em = 4.1E7 af = 1
+ ef = 0.84 kf = 0 lintnoi = -1E-7
+ tnoia = 1.5E7 tnoib = 9.9E6 ntnoi = 1
+ rnoia = 0.94 rnoib = 0.26 xpart = 0
+ cgso = {2.449068E-10/sw_func_tox_lv_ratio} cgdo = {2.449068E-10/sw_func_tox_lv_ratio} cgbo = {1E-13/sw_func_tox_lv_ratio}
+ ckappas = 0.6 cf = 1.4067E-12 clc = 1E-7
+ cle = 0.6 dlc = 9.87908E-9 dwc = 0
+ vfbcv = -1 noff = 3.4037 voffcv = -0.17287
+ acde = 0.4 moin = 6.9 cgsl = {0/sw_func_tox_lv_ratio}
+ cgdl = {0/sw_func_tox_lv_ratio} ijthsrev = 0.1 ijthsfwd = 0.1
+ xjbvs = 1 bvs = 11.7 jss = 2.75E-3
+ jsws = 6E-10 cjs = {sw_nsd_pw_cj} mjs = 0.44
+ mjsws = 9E-4 cjsws = {3.67354204E-11*sw_func_nsd_pw_cj} cjswgs = {2.38232788E-10*sw_func_nsd_pw_cj}
+ mjswgs = 0.8 pbs = 0.729 pbsws = 0.2
+ pbswgs = 0.95578 xrcrg1 = 12 xrcrg2 = 1
+ rbpb = 50 rbpd = 50 rbps = 50
+ rbdb = 50 rbsb = 50 gbmin = 1E-12
+ tnom = 30 ute = -2.03279478266222 lute = -2.15290845296312E-7
+ wute = 2.794027037788099E-7 pute = 2.696841465569178E-12 kt1 = -0.324283365527323
+ lkt1 = -2.448678831857541E-8 wkt1 = 2.731866969755221E-8 pkt1 = 3.104285936316088E-14
+ kt1l = 0 kt2 = -0.051806652019034 lkt2 = -2.455802143053303E-9
+ wkt2 = 2.691404929408572E-8 pkt2 = 1.361773604938209E-14 ua1 = 3.655919032718215E-10
+ lua1 = -2.536140922103683E-15 wua1 = -9.941278708174984E-16 pua1 = 1.052221902667555E-20
+ ub1 = -8.264202059134739E-19 lub1 = 3.027377223433322E-24 wub1 = 1.572841592195014E-24
+ pub1 = -9.612168782898868E-30 uc1 = 1.736274370701889E-11 luc1 = 1.253009184854528E-16
+ wuc1 = -2.281242334128314E-17 puc1 = -1.646606722397191E-22 at = 1.627603934958068E5
+ lat = -0.090498419952843 wat = 5.446948710511679E-3 pat = -2.165780885801907E-8
+ prt = 0 njs = 1.2928 xtis = 2
+ tpb = 1.2287E-3 tpbsw = 0 tpbswg = 0
+ tcj = 7.92E-4 tcjsw = 1E-5 tcjswg = 0
+ tvoff = 0 tvfbsdoff = 0 saref = 3E-6
+ sbref = 3E-6 wlod = 0 ku0 = -2.7E-8
+ kvsat = 0.2 kvth0 = 9.8E-9 tku0 = 0
+ llodku0 = 0 wlodku0 = 1 llodvth = 0
+ wlodvth = 1 lku0 = 0 wku0 = 0
+ pku0 = 0 lkvth0 = 0 wkvth0 = 2E-7
+ pkvth0 = 0 stk2 = 0 lodk2 = 1
+ steta0 = 0 lodeta0 = 1

.model nshort_model.28 nmos
+ level = 54 lmin = 1E-6 lmax = 2E-6 wmin = 1E-6
+ wmax = 3E-6 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 4.148E-9
+ toxm = 4.148E-9 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 9.999999999999999E22 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {2.1859E-8+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {1.1932E-8-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = 0 dwb = 0 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = 0.477523650628441 lvth0 = 8.962049081966782E-8
+ wvth0 = 4.72786256095353E-8 pvth0 = -3.318630002067166E-14 k1 = 0.645606612277521
+ lk1 = -1.230030867818668E-7 wk1 = -4.539006469691117E-8 pk1 = 6.661336302019187E-15
+ k2 = -0.063869778060352 lk2 = 3.953293735627536E-8 wk2 = 1.286178862136436E-8
+ pk2 = -3.774192821767429E-15 k3 = 2 k3b = 0.54
+ w0 = 0 lpe0 = 1.0325E-7 lpeb = -7.082E-8
+ vbm = -3 dvtp0 = 0 dvtp1 = 0
+ dvt0 = 0 dvt1 = 0.53 dvt2 = -0.032
+ dvt0w = -3.58 dvt1w = 1.6706E6 dvt2w = 0.068
+ vfbsdoff = 0 u0 = 0.035926649772123 lu0 = -1.016882188783929E-8
+ wu0 = -7.008272852595971E-9 pu0 = 5.903347369083766E-15 ua = 2.575128210417254E-10
+ lua = -1.738533746339784E-15 wua = -1.133298760196708E-15 pua = 1.229916987630127E-21
+ ub = 4.777618285137964E-19 lub = 1.804398229704163E-24 wub = 1.245483265139841E-24
+ pub = -1.435304544747932E-30 uc = 6.085907053182832E-11 luc = 1.588811313356571E-17
+ wuc = -2.145136882426745E-17 puc = 1.441305896009977E-23 ud = 0
+ up = 0 lp = 1 eu = 1.67
+ vsat = 9.103756266138205E4 lvsat = -0.021811724927413 wvsat = -0.019889635360472
+ pvsat = 3.930462446270118E-8 a0 = 2.441633676557941 la0 = -1.322191386157056E-6
+ wa0 = -9.809426784684994E-7 pa0 = 5.516662393195666E-13 ags = 0.064500372889099
+ lags = 1.312834779915688E-6 wags = 2.51193525481592E-7 pags = -9.333210958036527E-13
+ b0 = 6.155439406464786E-24 lb0 = -6.00854600046891E-30 wb0 = -5.886335906492957E-30
+ pb0 = 5.745864386420409E-36 b1 = 0 keta = 0.087985438064787
+ lketa = -1.643788790090274E-7 wketa = -1.097549215350126E-7 pketa = 1.911021403550948E-13
+ a1 = 0 a2 = 0.42385546 rdsw = 65.968
+ rdswmin = 0 rdw = 0 rdwmin = 0
+ rsw = 0 rswmin = 0 prwb = 0
+ prwg = 0.021507 wr = 1 voff = -0.053511380065817
+ lvoff = -7.014845472138018E-8 wvoff = -4.537880931830508E-8 pvoff = 2.005836458480078E-14
+ voffl = 5.8197729E-9 minv = 0 nfactor = 3.489757690952624
+ lnfactor = -9.275576208690838E-7 wnfactor = -6.428656023039206E-7 pnfactor = 8.400364844236369E-14
+ eta0 = 0.155620059086532 leta0 = -1.494355210830233E-7 peta0 = 1.36332377606075E-19
+ etab = -0.055968045 letab = -2.772905142588E-8 dsub = 0.8528408
+ ldsub = -5.786932471488001E-7 cit = 0 cdsc = 0
+ cdscb = 0 cdscd = 5.4E-3 pclm = -0.015785938518114
+ lpclm = 9.771797303218076E-7 wpclm = 4.253421582428692E-7 ppclm = -6.924048793658232E-13
+ pdiblc1 = 0.033377126812219 lpdiblc1 = 7.047352981298092E-7 wpdiblc1 = 3.889142858164725E-7
+ ppdiblc1 = -7.685475211162206E-13 pdiblc2 = 7.136341112324988E-3 lpdiblc2 = -4.943605032876209E-9
+ wpdiblc2 = -2.234852584056031E-9 ppdiblc2 = 5.667812464254645E-15 pdiblcb = -0.072170518049902
+ lpdiblcb = 9.321535885706112E-8 wpdiblcb = 6.785913988186195E-8 ppdiblcb = -1.340988892495831E-13
+ drout = 0.916922828629243 ldrout = -7.053280508760772E-7 wdrout = -1.894445477601146E-7
+ pdrout = 3.743681908324818E-13 pscbe1 = 1.324356440665688E9 lpscbe1 = -1.060556841194948E3
+ wpscbe1 = -501.432625792666 ppscbe1 = 1.014191417211587E-3 pscbe2 = 1E-12
+ pvag = 0 delta = 0.01 fprout = 0
+ pdits = 0 pditsl = 0 pditsd = 0
+ lambda = 0 vtl = 0 lc = 5E-9
+ xn = 3 alpha0 = -1.211463609528001E-8 lalpha0 = 8.322424851478224E-14
+ walpha0 = 4.139362197808895E-14 palpha0 = -8.179942656129277E-20 alpha1 = 0.459716683452176
+ lalpha1 = 7.712529120295508E-7 walpha1 = 5.160404873268423E-7 palpha1 = -1.019766184464117E-12
+ beta0 = 12.894722215715255 lbeta0 = 1.907520179525318E-6 wbeta0 = 9.230777701113843E-7
+ pbeta0 = -1.82412721231683E-12 aigbacc = 1 bigbacc = 0
+ cigbacc = 0 nigbacc = 0 aigbinv = 0.35
+ bigbinv = 0.03 cigbinv = 6E-3 eigbinv = 1.1
+ nigbinv = 0 aigc = 0.43 bigc = 0.054
+ cigc = 0.075 aigsd = 0.43 bigsd = 0.054
+ cigsd = 0.075 dlcig = 0 nigc = 0
+ poxedge = 1 pigcd = 1 ntox = 1
+ toxref = 4.148E-9 agidl = 0 bgidl = 2.3E9
+ cgidl = 0.5 egidl = 0.8 noia = 2.5E42
+ noib = 0 noic = 0 em = 4.1E7
+ af = 1 ef = 0.84 kf = 0
+ lintnoi = -1E-7 tnoia = 1.5E7 tnoib = 9.9E6
+ ntnoi = 1 rnoia = 0.94 rnoib = 0.26
+ xpart = 0 cgso = {2.449068E-10/sw_func_tox_lv_ratio} cgdo = {2.449068E-10/sw_func_tox_lv_ratio}
+ cgbo = {1E-13/sw_func_tox_lv_ratio} ckappas = 0.6 cf = 1.4067E-12
+ clc = 1E-7 cle = 0.6 dlc = 9.87908E-9
+ dwc = 0 vfbcv = -1 noff = 3.4037
+ voffcv = -0.17287 acde = 0.4 moin = 6.9
+ cgsl = {0/sw_func_tox_lv_ratio} cgdl = {0/sw_func_tox_lv_ratio} ijthsrev = 0.1
+ ijthsfwd = 0.1 xjbvs = 1 bvs = 11.7
+ jss = 2.75E-3 jsws = 6E-10 cjs = {sw_nsd_pw_cj}
+ mjs = 0.44 mjsws = 9E-4 cjsws = {3.67354204E-11*sw_func_nsd_pw_cj}
+ cjswgs = {2.38232788E-10*sw_func_nsd_pw_cj} mjswgs = 0.8 pbs = 0.729
+ pbsws = 0.2 pbswgs = 0.95578 xrcrg1 = 12
+ xrcrg2 = 1 rbpb = 50 rbpd = 50
+ rbps = 50 rbdb = 50 rbsb = 50
+ gbmin = 1E-12 tnom = 30 ute = -3.0277394274369
+ lute = 1.750855085250148E-6 wute = 3.074160143516359E-6 pute = -2.825979322364022E-12
+ kt1 = -0.417237722725245 lkt1 = 1.592036632970971E-7 wkt1 = 8.736010672936857E-8
+ pkt1 = -8.760718584714455E-14 kt1l = 0 kt2 = -0.070041060074391
+ lkt2 = 3.357786805382801E-8 wkt2 = 6.734918641351626E-8 pkt2 = -6.628759407726089E-14
+ ua1 = -3.589986593100069E-9 lua1 = 5.280620145402677E-15 wua1 = 9.092962842073589E-15
+ pua1 = -9.411244066334185E-21 ub1 = 3.126782379401146E-18 lub1 = -4.78468872069997E-24
+ wub1 = -7.444164388696672E-24 pub1 = 8.206661348156504E-30 uc1 = 1.899569500110689E-10
+ luc1 = -2.157687059834073E-16 wuc1 = -2.556053943821315E-16 puc1 = 2.953698983810588E-22
+ at = 1.764487322965764E5 lat = -0.117548439037241 wat = -0.038606927335354
+ pat = 6.539864153575358E-8 prt = 0 njs = 1.2928
+ xtis = 2 tpb = 1.2287E-3 tpbsw = 0
+ tpbswg = 0 tcj = 7.92E-4 tcjsw = 1E-5
+ tcjswg = 0 tvoff = 0 tvfbsdoff = 0
+ saref = 3E-6 sbref = 3E-6 wlod = 0
+ ku0 = -2.7E-8 kvsat = 0.2 kvth0 = 9.8E-9
+ tku0 = 0 llodku0 = 0 wlodku0 = 1
+ llodvth = 0 wlodvth = 1 lku0 = 0
+ wku0 = 0 pku0 = 0 lkvth0 = 0
+ wkvth0 = 2E-7 pkvth0 = 0 stk2 = 0
+ lodk2 = 1 steta0 = 0 lodeta0 = 1

.model nshort_model.29 nmos
+ level = 54 lmin = 5E-7 lmax = 1E-6 wmin = 1E-6
+ wmax = 3E-6 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 4.148E-9
+ toxm = 4.148E-9 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 9.999999999999999E22 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {2.1859E-8+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {1.1932E-8-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = 0 dwb = 0 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = 0.566059628514088 lvth0 = 3.197335510283302E-9
+ wvth0 = 2.003032891864236E-8 pvth0 = -6.588256682010195E-15 k1 = 0.458516519101106
+ lk1 = 5.962228841098677E-8 wk1 = -5.685125468342146E-8 pk1 = 1.78490164506914E-14
+ k2 = -4.145550992556365E-3 lk2 = -1.876603075677392E-8 wk2 = 1.024776896284332E-8
+ pk2 = -1.222554128377333E-15 k3 = 2 k3b = 0.54
+ w0 = 0 lpe0 = 1.0325E-7 lpeb = -7.082E-8
+ vbm = -3 dvtp0 = 0 dvtp1 = 0
+ dvt0 = 0 dvt1 = 0.53 dvt2 = -0.032
+ dvt0w = -3.58 dvt1w = 1.6706E6 dvt2w = 0.068
+ vfbsdoff = 0 u0 = 0.027990003623927 lu0 = -2.421575863324163E-9
+ wu0 = -1.087917847751013E-9 pu0 = 1.242757160744279E-16 ua = -1.40570005382719E-9
+ lua = -1.150117835167402E-16 wua = 1.001024272548275E-16 pua = 2.594968611593532E-23
+ ub = 2.338303153681471E-18 lub = -1.174313727971054E-26 wub = -1.18860460318465E-25
+ pub = -1.035195179539629E-31 uc = 7.919268734926569E-11 luc = -2.007990252140323E-18
+ wuc = -1.538819451144927E-17 puc = 8.494576239082681E-24 ud = 0
+ up = 0 lp = 1 eu = 1.67
+ vsat = 1.2948289910273E4 lvsat = 0.054414025418764 wvsat = 0.042173633651607
+ pvsat = -2.127756669767319E-8 a0 = 0.693942288687013 la0 = 3.837930944337201E-7
+ wa0 = -8.117344461399211E-7 pa0 = 3.864959922472775E-13 ags = 1.583106305469726
+ lags = -1.695311406898341E-7 wags = -1.256175984351775E-6 pags = 5.380765480470508E-13
+ b0 = 0 b1 = 0 keta = -0.121329301874515
+ lketa = 3.994077397636312E-8 wketa = 1.626512554193175E-7 pketa = -7.480333559239716E-14
+ a1 = 0 a2 = 0.42385546 rdsw = 65.968
+ rdswmin = 0 rdw = 0 rdwmin = 0
+ rsw = 0 rswmin = 0 prwb = 0
+ prwg = 0.021507 wr = 1 voff = -0.114730037551805
+ lvoff = -1.039071927763831E-8 wvoff = -4.038236408492458E-8 pvoff = 1.518115452046967E-14
+ voffl = 5.8197729E-9 minv = 0 nfactor = 2.436604371838811
+ lnfactor = 1.004632474373957E-7 wnfactor = -1.52331479270948E-6 pnfactor = 9.434417993680858E-13
+ eta0 = -0.461671638173064 leta0 = 4.5312512711317E-7 peta0 = -6.569664531404419E-20
+ etab = -0.163985492410515 letab = 7.771066761963047E-8 wetab = -4.206422396178857E-10
+ petab = 4.106040332116445E-16 dsub = 0.185943845767231 ldsub = 7.228887816815831E-8
+ wdsub = 2.223041067201484E-8 pdsub = -2.169990415173788E-14 cit = 0
+ cdsc = 0 cdscb = 0 cdscd = 5.4E-3
+ pclm = 1.58816424351618 lpclm = -5.884937845684198E-7 wpclm = -6.890316894522496E-7
+ ppclm = 3.953755508278994E-13 pdiblc1 = 0.835545369741637 lpdiblc1 = -7.829000185034106E-8
+ wpdiblc1 = -2.961010697942895E-7 ppdiblc1 = -9.987937195175382E-14 pdiblc2 = 3.236684340266956E-3
+ lpdiblc2 = -1.13700967002657E-9 wpdiblc2 = 6.283115830305821E-9 ppdiblc2 = -2.646883151866876E-15
+ pdiblcb = 0.069341036099804 lpdiblcb = -4.491916356441626E-8 wpdiblcb = -1.357182797637238E-7
+ ppdiblcb = 6.462035885358042E-14 drout = -0.572845337258485 ldrout = 7.488882875009059E-7
+ wdrout = 3.78889095520229E-7 pdrout = -1.804027383846197E-13 pscbe1 = -2.974272852586101E8
+ lpscbe1 = 522.5246378938936 wpscbe1 = 1.049449959201674E3 ppscbe1 = -4.996809057744484E-4
+ pscbe2 = 1E-12 pvag = 0 delta = 0.01
+ fprout = 0 pdits = 0 pditsl = 0
+ pditsd = 0 lambda = 0 vtl = 0
+ lc = 5E-9 xn = 3 alpha0 = -4.404141966999357E-6
+ lalpha0 = 4.370440239194166E-12 walpha0 = 4.238049841398835E-12 palpha0 = -4.178306641961782E-18
+ alpha1 = 1.630566633095648 lalpha1 = -3.716558744156293E-7 walpha1 = -1.032080974653684E-6
+ palpha1 = 4.914109069477066E-13 beta0 = 9.937786841917873 lbeta0 = 4.7938912475624E-6
+ wbeta0 = 3.750741843237092E-6 pbeta0 = -4.584311910001466E-12 aigbacc = 1
+ bigbacc = 0 cigbacc = 0 nigbacc = 0
+ aigbinv = 0.35 bigbinv = 0.03 cigbinv = 6E-3
+ eigbinv = 1.1 nigbinv = 0 aigc = 0.43
+ bigc = 0.054 cigc = 0.075 aigsd = 0.43
+ bigsd = 0.054 cigsd = 0.075 dlcig = 0
+ nigc = 0 poxedge = 1 pigcd = 1
+ ntox = 1 toxref = 4.148E-9 agidl = 0
+ bgidl = 2.3E9 cgidl = 0.5 egidl = 0.8
+ noia = 2.5E42 noib = 0 noic = 0
+ em = 4.1E7 af = 1 ef = 0.84
+ kf = 0 lintnoi = -1E-7 tnoia = 1.5E7
+ tnoib = 9.9E6 ntnoi = 1 rnoia = 0.94
+ rnoib = 0.26 xpart = 0 cgso = {2.449068E-10/sw_func_tox_lv_ratio}
+ cgdo = {2.449068E-10/sw_func_tox_lv_ratio} cgbo = {1E-13/sw_func_tox_lv_ratio} ckappas = 0.6
+ cf = 1.4067E-12 clc = 1E-7 cle = 0.6
+ dlc = 9.87908E-9 dwc = 0 vfbcv = -1
+ noff = 3.4037 voffcv = -0.17287 acde = 0.4
+ moin = 6.9 cgsl = {0/sw_func_tox_lv_ratio} cgdl = {0/sw_func_tox_lv_ratio}
+ ijthsrev = 0.1 ijthsfwd = 0.1 xjbvs = 1
+ bvs = 11.7 jss = 2.75E-3 jsws = 6E-10
+ cjs = {sw_nsd_pw_cj} mjs = 0.44 mjsws = 9E-4
+ cjsws = {3.67354204E-11*sw_func_nsd_pw_cj} cjswgs = {2.38232788E-10*sw_func_nsd_pw_cj} mjswgs = 0.8
+ pbs = 0.729 pbsws = 0.2 pbswgs = 0.95578
+ xrcrg1 = 12 xrcrg2 = 1 rbpb = 50
+ rbpd = 50 rbps = 50 rbdb = 50
+ rbsb = 50 gbmin = 1E-12 tnom = 30
+ ute = -1.203670483319997 lute = -2.968427758435071E-8 wute = 3.131493981194432E-7
+ pute = -1.308573373952585E-13 kt1 = -0.226461056862881 lkt1 = -2.702030821112777E-8
+ wkt1 = -1.599906771944424E-8 pkt1 = 1.328542526262179E-14 kt1l = 0
+ kt2 = -0.034162380533053 lkt2 = -1.444602678935926E-9 wkt2 = -1.86181061502071E-9
+ pkt2 = 1.271751718187074E-15 ua1 = 2.584303227153219E-9 lua1 = -7.463264225800863E-16
+ wua1 = -1.140466426648708E-15 pua1 = 5.779746463193232E-22 ub1 = -2.95942821024612E-18
+ lub1 = 1.156280539435955E-24 wub1 = 2.015772679931911E-24 pub1 = -1.027523782266326E-30
+ uc1 = -1.160809765777988E-10 luc1 = 8.296593152534369E-17 wuc1 = 1.089993776735146E-16
+ puc1 = -6.053394539425141E-23 at = 6.661975032709845E4 lat = -0.010340415893483
+ wat = 0.050665234998831 pat = -2.17431299164886E-8 prt = 0
+ njs = 1.2928 xtis = 2 tpb = 1.2287E-3
+ tpbsw = 0 tpbswg = 0 tcj = 7.92E-4
+ tcjsw = 1E-5 tcjswg = 0 tvoff = 0
+ tvfbsdoff = 0 saref = 2.75E-6 sbref = 2.74E-6
+ wlod = 0 ku0 = -2.7E-8 kvsat = 0.2
+ kvth0 = 9.8E-9 tku0 = 0 llodku0 = 0
+ wlodku0 = 1 llodvth = 0 wlodvth = 1
+ lku0 = 0 wku0 = 0 pku0 = 0
+ lkvth0 = 0 wkvth0 = 2E-7 pkvth0 = 0
+ stk2 = 0 lodk2 = 1 steta0 = 0
+ lodeta0 = 1

.model nshort_model.30 nmos
+ level = 54 lmin = 2.5E-7 lmax = 5E-7 wmin = 1E-6
+ wmax = 3E-6 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 4.148E-9
+ toxm = 4.148E-9 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 9.999999999999999E22 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {2.1859E-8+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {1.1932E-8-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = 0 dwb = 0 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = 0.612651989599055 lvth0 = -1.898696492726835E-8
+ wvth0 = 8.028887824505228E-9 pvth0 = -8.739385252121171E-16 k1 = 0.462637129932164
+ lk1 = 5.766031725232988E-8 wk1 = -2.007586278331666E-7 pk1 = 8.636849747271844E-14
+ k2 = -0.021752529221711 lk2 = -1.038271457065718E-8 wk2 = 7.696065741008098E-8
+ pk2 = -3.298696198209128E-14 k3 = 2 k3b = 0.54
+ w0 = 0 lpe0 = 1.0325E-7 lpeb = -7.082E-8
+ vbm = -3 dvtp0 = 0 dvtp1 = 0
+ dvt0 = 0 dvt1 = 0.53 dvt2 = -0.032
+ dvt0w = -3.58 dvt1w = 1.6706E6 dvt2w = 0.068
+ vfbsdoff = 0 u0 = 0.032295809074906 lu0 = -4.471724847531677E-9
+ wu0 = -1.236184285987223E-8 pu0 = 5.492197275645774E-15 ua = -8.479286303324799E-10
+ lua = -3.805868380138177E-16 wua = -8.799753120629196E-16 pua = 4.925999806037301E-22
+ ub = 1.912286419330101E-18 lub = 1.910987665474136E-25 wub = 1.966556271993666E-25
+ pub = -2.537480858003531E-31 uc = 8.333407064379076E-11 luc = -3.979851928462318E-18
+ wuc = -1.853305262741369E-17 puc = 9.991956402985515E-24 ud = 0
+ up = 0 lp = 1 eu = 1.67
+ vsat = 1.111055746967808E5 lvsat = 7.677808469655045E-3 wvsat = -0.019250865289302
+ pvsat = 7.968848530055419E-9 a0 = 1.5 ags = 2.851481720546714
+ lags = -7.734503373229315E-7 wags = -1.813402463997012E-6 pags = 8.033921351594153E-13
+ b0 = 0 b1 = 0 keta = -0.053901431379012
+ lketa = 7.835937430116379E-9 wketa = 6.583485076519725E-8 pketa = -2.870555994600298E-14
+ a1 = 0 a2 = 0.42385546 rdsw = 65.968
+ rdswmin = 0 rdw = 0 rdwmin = 0
+ rsw = 0 rswmin = 0 prwb = 0
+ prwg = 0.021507 wr = 1 voff = -0.143325501560755
+ lvoff = 3.224610573727276E-9 wvoff = 2.655778815997409E-8 pvoff = -1.66914618088074E-14
+ voffl = 5.8197729E-9 minv = 0 nfactor = 1.997280892146944
+ lnfactor = 3.096409717639626E-7 wnfactor = 1.782742242576902E-6 pnfactor = -6.306909731850309E-13
+ eta0 = 0.278375424628437 leta0 = 1.007620788191146E-7 weta0 = 6.256219229285958E-7
+ peta0 = -2.978811198955298E-13 etab = -0.019668379145861 letab = 8.996094578250979E-9
+ wetab = 5.629759898808305E-8 petab = -2.659499247198096E-14 dsub = 0.074886354620701
+ ldsub = 1.251673477727024E-7 wdsub = 1.023823799982279E-7 pdsub = -5.986314221884363E-14
+ cit = 0 cdsc = 0 cdscb = 0
+ cdscd = 3.951991430587008E-3 lcdscd = 6.894490082060244E-10 wcdscd = 4.280721669601379E-9
+ pcdscd = -2.038205692877322E-15 pclm = 0.344302754572617 lpclm = 3.753449331212422E-9
+ wpclm = 3.750271998358021E-7 ppclm = -1.112611924821563E-13 pdiblc1 = 1.224782807096824
+ lpdiblc1 = -2.636199583228907E-7 wpdiblc1 = -1.221179610852325E-6 ppdiblc1 = 3.405838242734549E-13
+ pdiblc2 = 1.800516138135236E-3 lpdiblc2 = -4.531982869363818E-10 wpdiblc2 = -6.068438370389481E-9
+ ppdiblc2 = 3.234136459035382E-15 pdiblcb = 0.208545827471269 lpdiblcb = -1.111995761088603E-7
+ wpdiblcb = -1.556098968468191E-7 ppdiblcb = 7.409147384505703E-14 drout = 0.785188992676532
+ ldrout = 1.02279253782967E-7 wdrout = 6.350419143522381E-7 pdrout = -3.023663169320172E-13
+ pscbe1 = 7.96289101766251E8 lpscbe1 = 1.766892241424334 wpscbe1 = 10.970461652264092
+ ppscbe1 = -5.223431729262415E-6 pscbe2 = 1E-12 pvag = 0
+ delta = 0.01 fprout = 0 pdits = 0
+ pditsl = 0 pditsd = 0 lambda = 0
+ vtl = 0 lc = 5E-9 xn = 3
+ alpha0 = 4.690976999227045E-6 lalpha0 = 3.992667509099126E-14 walpha0 = -4.44994241395341E-12
+ palpha0 = -4.164076146738636E-20 alpha1 = 0.85 beta0 = 18.722278759315106
+ lbeta0 = 6.112784039805503E-7 wbeta0 = -5.04760926340305E-6 pbeta0 = -3.951002074902558E-13
+ aigbacc = 1 bigbacc = 0 cigbacc = 0
+ nigbacc = 0 aigbinv = 0.35 bigbinv = 0.03
+ cigbinv = 6E-3 eigbinv = 1.1 nigbinv = 0
+ aigc = 0.43 bigc = 0.054 cigc = 0.075
+ aigsd = 0.43 bigsd = 0.054 cigsd = 0.075
+ dlcig = 0 nigc = 0 poxedge = 1
+ pigcd = 1 ntox = 1 toxref = 4.148E-9
+ agidl = 0 bgidl = 2.3E9 cgidl = 0.5
+ egidl = 0.8 noia = 2.5E42 noib = 0
+ noic = 0 em = 4.1E7 af = 1
+ ef = 0.84 kf = 0 lintnoi = -1E-7
+ tnoia = 1.5E7 tnoib = 9.9E6 ntnoi = 1
+ rnoia = 0.94 rnoib = 0.26 xpart = 0
+ cgso = {2.449068E-10/sw_func_tox_lv_ratio} cgdo = {2.449068E-10/sw_func_tox_lv_ratio} cgbo = {1E-13/sw_func_tox_lv_ratio}
+ ckappas = 0.6 cf = 1.4067E-12 clc = 1E-7
+ cle = 0.6 dlc = 9.87908E-9 dwc = 0
+ vfbcv = -1 noff = 3.4037 voffcv = -0.17287
+ acde = 0.4 moin = 6.9 cgsl = {0/sw_func_tox_lv_ratio}
+ cgdl = {0/sw_func_tox_lv_ratio} ijthsrev = 0.1 ijthsfwd = 0.1
+ xjbvs = 1 bvs = 11.7 jss = 2.75E-3
+ jsws = 6E-10 cjs = {sw_nsd_pw_cj} mjs = 0.44
+ mjsws = 9E-4 cjsws = {3.67354204E-11*sw_func_nsd_pw_cj} cjswgs = {2.38232788E-10*sw_func_nsd_pw_cj}
+ mjswgs = 0.8 pbs = 0.729 pbsws = 0.2
+ pbswgs = 0.95578 xrcrg1 = 12 xrcrg2 = 1
+ rbpb = 50 rbpd = 50 rbps = 50
+ rbdb = 50 rbsb = 50 gbmin = 1E-12
+ tnom = 30 ute = -2.606566067562492 lute = 6.382848143145335E-7
+ wute = 1.400792392785474E-6 pute = -6.487233223035635E-13 kt1 = -0.314259011657515
+ lkt1 = 1.478345879297011E-8 wkt1 = 1.581645244202854E-8 pkt1 = -1.86308924498121E-15
+ kt1l = 0 kt2 = -0.06045385097825 lkt2 = 1.107371289295872E-8
+ wkt2 = 1.658720401007224E-8 pkt2 = -7.51248830934618E-15 ua1 = -1.266999316812888E-9
+ lua1 = 1.08741736549376E-15 wua1 = 3.224015306623059E-15 pua1 = -1.500112228233763E-21
+ ub1 = 1.225820583340563E-18 lub1 = -8.364670801472342E-25 wub1 = -3.022433145683173E-24
+ pub1 = 1.371347386718738E-30 uc1 = 1.065646913553946E-10 luc1 = -2.304368622169525E-17
+ wuc1 = -1.578243337277248E-16 puc1 = 6.651042925748913E-23 at = 6.75994436198608E4
+ lat = -0.010806883139125 wat = 1.814202621998158E-3 pat = 1.516605235287198E-9
+ prt = 0 njs = 1.2928 xtis = 2
+ tpb = 1.2287E-3 tpbsw = 0 tpbswg = 0
+ tcj = 7.92E-4 tcjsw = 1E-5 tcjswg = 0
+ tvoff = 0 tvfbsdoff = 0 saref = 1.75E-6
+ sbref = 1.74E-6 wlod = 0 ku0 = -2.7E-8
+ kvsat = 0.2 kvth0 = 9.8E-9 tku0 = 0
+ llodku0 = 0 wlodku0 = 1 llodvth = 0
+ wlodvth = 1 lku0 = 0 wku0 = 0
+ pku0 = 0 lkvth0 = 0 wkvth0 = 2E-7
+ pkvth0 = 0 stk2 = 0 lodk2 = 1
+ steta0 = 0 lodeta0 = 1

.model nshort_model.31 nmos
+ level = 54 lmin = 1.8E-7 lmax = 2.5E-7 wmin = 1E-6
+ wmax = 3E-6 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 4.148E-9
+ toxm = 4.148E-9 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 9.999999999999999E22 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {2.1859E-8+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {1.1932E-8-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = 0 dwb = 0 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = 0.619169315967313 lvth0 = -2.04607670428808E-8
+ wvth0 = -2.016353461842927E-9 pvth0 = 1.397652158317509E-15 k1 = 0.295034297600426
+ lk1 = 9.556135134449995E-8 wk1 = 5.852820629862499E-7 pk1 = -9.13836001864211E-14
+ k2 = 0.071441784150712 lk2 = -3.145730381944343E-8 wk2 = -2.18414505177594E-7
+ pk2 = 3.38079957848352E-14 k3 = 2 k3b = 0.54
+ w0 = 0 lpe0 = 1.0325E-7 lpeb = -7.082E-8
+ vbm = -3 dvtp0 = 0 dvtp1 = 0
+ dvt0 = 0 dvt1 = 0.53 dvt2 = -0.032
+ dvt0w = -3.58 dvt1w = 1.6706E6 dvt2w = 0.068
+ vfbsdoff = 0 u0 = -0.024636365367997 lu0 = 8.402689352288705E-9
+ wu0 = 4.475430299493788E-8 pu0 = -7.423819483377563E-15 ua = -5.524865571507865E-9
+ lua = 6.770369741158192E-16 wua = 4.171320034745794E-15 pua = -6.496797439422053E-22
+ ub = 3.885210836450437E-18 lub = -2.550504694425107E-25 wub = -2.31089753071306E-24
+ pub = 3.132999551173314E-31 uc = 1.329141934413475E-10 luc = -1.519170257741061E-17
+ wuc = -7.619479048656099E-17 puc = 2.303135115550165E-23 ud = 0
+ up = 0 lp = 1 eu = 1.67
+ vsat = 1.583898243529192E5 lvsat = -3.014862610585462E-3 wvsat = -0.031785628970978
+ pvsat = 1.080340984997489E-8 a0 = 1.5 ags = -4.62568095664828
+ lags = 9.174053218472357E-7 wags = 5.61880793658553E-6 pags = -8.772981959867183E-13
+ b0 = 0 b1 = 0 keta = 0.063506330926503
+ lketa = -1.871418430660354E-8 wketa = -2.344106101206024E-7 pketa = 3.919074759686821E-14
+ a1 = 0 a2 = 0.42385546 rdsw = 65.968
+ rdswmin = 0 rdw = 0 rdwmin = 0
+ rsw = 0 rswmin = 0 prwb = 0
+ prwg = 0.021507 wr = 1 voff = -0.03809148782817
+ lvoff = -2.057258835570468E-8 wvoff = -7.228733796062234E-8 pvoff = 5.660979631599795E-15
+ voffl = 5.8197729E-9 minv = 0 nfactor = 4.242082229265567
+ lnfactor = -1.979894234066945E-7 wnfactor = 3.777650498068708E-7 pnfactor = -3.129750507207872E-13
+ eta0 = 2.337205764411024 leta0 = -3.648135788979605E-7 weta0 = -2.234364006612762E-6
+ peta0 = 3.488646582672346E-13 etab = 0.186731340267605 letab = -3.767831237103244E-8
+ wetab = -2.206423149697856E-7 petab = 3.603109191079563E-14 dsub = 1.007040371219926
+ ldsub = -8.562623292497989E-8 wdsub = -5.244244295876621E-7 pdsub = 8.188044247367117E-14
+ cit = 0 cdsc = 0 cdscb = 0
+ cdscd = 0.01491365114832 lcdscd = -1.789376873723244E-9 wcdscd = -1.229936548341775E-8
+ pcdscd = 1.711148895557811E-15 pclm = 0.462351362810255 lpclm = -2.294159074121403E-8
+ wpclm = 1.830701292617419E-8 ppclm = -3.05939162951607E-14 pdiblc1 = -0.605552529566332
+ lpdiblc1 = 1.502847533687688E-7 wpdiblc1 = 9.20445025625051E-7 ppdiblc1 = -1.43714604520993E-13
+ pdiblc2 = -0.019407621262409 lpdiblc2 = 4.342725072273097E-9 wpdiblc2 = 2.659777256727123E-8
+ ppdiblc2 = -4.152869817563462E-15 pdiblcb = -0.684452407472819 lpdiblcb = 9.073947274845608E-8
+ wpdiblcb = 5.557496315957824E-7 ppdiblcb = -8.677252447883908E-14 drout = 2.875019149215816
+ ldrout = -3.703065784962007E-7 wdrout = -2.268006836972279E-6 pdrout = 3.541175154975038E-13
+ pscbe1 = 8.32391288210818E8 lpscbe1 = -6.397111792404282 wpscbe1 = -39.18022018665748
+ ppscbe1 = 6.117442859063952E-6 pscbe2 = 1E-12 pvag = 0
+ delta = 0.01 fprout = 0 pdits = 0
+ pditsl = 0 pditsd = 0 lambda = 0
+ vtl = 0 lc = 5E-9 xn = 3
+ alpha0 = 1.5648775251336E-5 lalpha0 = -2.43802599044792E-12 walpha0 = -1.49439864036981E-11
+ palpha0 = 2.331440370197517E-18 alpha1 = 0.85 beta0 = 37.249003993673035
+ lbeta0 = -3.578281133616213E-6 wbeta0 = -2.141467363815649E-5 pbeta0 = 3.306082261958987E-12
+ aigbacc = 1 bigbacc = 0 cigbacc = 0
+ nigbacc = 0 aigbinv = 0.35 bigbinv = 0.03
+ cigbinv = 6E-3 eigbinv = 1.1 nigbinv = 0
+ aigc = 0.43 bigc = 0.054 cigc = 0.075
+ aigsd = 0.43 bigsd = 0.054 cigsd = 0.075
+ dlcig = 0 nigc = 0 poxedge = 1
+ pigcd = 1 ntox = 1 toxref = 4.148E-9
+ agidl = 0 bgidl = 2.3E9 cgidl = 0.5
+ egidl = 0.8 noia = 2.5E42 noib = 0
+ noic = 0 em = 4.1E7 af = 1
+ ef = 0.84 kf = 0 lintnoi = -1E-7
+ tnoia = 1.5E7 tnoib = 9.9E6 ntnoi = 1
+ rnoia = 0.94 rnoib = 0.26 xpart = 0
+ cgso = {2.449068E-10/sw_func_tox_lv_ratio} cgdo = {2.449068E-10/sw_func_tox_lv_ratio} cgbo = {1E-13/sw_func_tox_lv_ratio}
+ ckappas = 0.6 cf = 1.4067E-12 clc = 1E-7
+ cle = 0.6 dlc = 9.87908E-9 dwc = 0
+ vfbcv = -1 noff = 3.4037 voffcv = -0.17287
+ acde = 0.4 moin = 6.9 cgsl = {0/sw_func_tox_lv_ratio}
+ cgdl = {0/sw_func_tox_lv_ratio} ijthsrev = 0.1 ijthsfwd = 0.1
+ xjbvs = 1 bvs = 11.7 jss = 2.75E-3
+ jsws = 6E-10 cjs = {sw_nsd_pw_cj} mjs = 0.44
+ mjsws = 9E-4 cjsws = {3.67354204E-11*sw_func_nsd_pw_cj} cjswgs = {2.38232788E-10*sw_func_nsd_pw_cj}
+ mjswgs = 0.8 pbs = 0.729 pbsws = 0.2
+ pbswgs = 0.95578 xrcrg1 = 12 xrcrg2 = 1
+ rbpb = 50 rbpd = 50 rbps = 50
+ rbdb = 50 rbsb = 50 gbmin = 1E-12
+ tnom = 30 ute = 3.639950273363172 lute = -7.742774049570323E-7
+ wute = -4.742196196694681E-6 pute = 7.404275453671207E-13 kt1 = -0.233589439068766
+ lkt1 = -3.458835673959137E-9 wkt1 = -7.049042397122212E-9 pkt1 = 3.307622295964991E-15
+ kt1l = 0 kt2 = 0.02731375525493 lkt2 = -8.773702510187703E-9
+ wkt2 = -5.373606204749268E-8 pkt2 = 8.390133783847316E-15 ua1 = 1.149466622343795E-8
+ lua1 = -1.798454633116404E-15 wua1 = -1.101494718364644E-14 pua1 = 1.719829793465821E-21
+ ub1 = -9.568152366629329E-18 lub1 = 1.604438786867156E-24 wub1 = 9.826663498378966E-24
+ pub1 = -1.534295931982898E-30 uc1 = -3.132377929621681E-10 luc1 = 7.188876837194107E-17
+ wuc1 = 4.40295224651948E-16 puc1 = -6.874593519625655E-23 at = -1.208962094653769E5
+ lat = 0.031818769866958 wat = 0.074819732539818 pat = -1.499257327820886E-8
+ prt = 0 njs = 1.2928 xtis = 2
+ tpb = 1.2287E-3 tpbsw = 0 tpbswg = 0
+ tcj = 7.92E-4 tcjsw = 1E-5 tcjswg = 0
+ tvoff = 0 tvfbsdoff = 0 saref = 1.25E-6
+ sbref = 1.24E-6 wlod = 0 ku0 = -2.7E-8
+ kvsat = 0.2 kvth0 = 9.8E-9 tku0 = 0
+ llodku0 = 0 wlodku0 = 1 llodvth = 0
+ wlodvth = 1 lku0 = 0 wku0 = 0
+ pku0 = 0 lkvth0 = 0 wkvth0 = 2E-7
+ pkvth0 = 0 stk2 = 0 lodk2 = 1
+ steta0 = 0 lodeta0 = 1

.model nshort_model.32 nmos
+ level = 54 lmin = 1.5E-7 lmax = 1.8E-7 wmin = 1E-6
+ wmax = 3E-6 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 4.148E-9
+ toxm = 4.148E-9 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 9.999999999999999E22 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {2.1859E-8+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {1.1932E-8-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = 0 dwb = 0 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = 0.759048887425729 lvth0 = -4.230100381211201E-8
+ wvth0 = -1.6256345045912E-7 pvth0 = 2.646483369508436E-14 k1 = 0.90707349
+ k2 = -0.126764169876655 lk2 = -5.102189814265024E-10 wk2 = -1.92983060643618E-8
+ pk2 = 2.718788920091567E-15 k3 = 2 k3b = 0.54
+ w0 = 0 lpe0 = 1.0325E-7 lpeb = -7.082E-8
+ vbm = -3 dvtp0 = 0 dvtp1 = 0
+ dvt0 = 0 dvt1 = 0.53 dvt2 = -0.032
+ dvt0w = -3.58 dvt1w = 1.6706E6 dvt2w = 0.068
+ vfbsdoff = 0 u0 = 0.041098529733864 lu0 = -1.860894229335405E-9
+ wu0 = -1.430479191079305E-8 pu0 = 1.797431358823641E-15 ua = -1.228006274061534E-9
+ lua = 6.1425508497389E-18 wua = 4.723924745508983E-17 pua = -5.762266137783807E-24
+ ub = 3.523075930692824E-18 lub = -1.985081737971401E-25 wub = -1.145501098600934E-24
+ pub = 1.313396177930725E-31 uc = -2.302186543625218E-11 luc = 9.155529911502298E-18
+ wuc = 2.446644567936146E-16 puc = -2.706632827783584E-23 ud = 0
+ up = 0 lp = 1 eu = 1.67
+ vsat = 5.599549984204079E4 lvsat = 0.012972577641245 wvsat = 0.105678660575932
+ pvsat = -1.065971446272146E-8 a0 = 1.5 ags = 1.25
+ b0 = 0 b1 = 0 keta = -0.407751228592621
+ lketa = 5.486608600647437E-8 wketa = 1.958221001234087E-7 pketa = -2.798406684979071E-14
+ a1 = 0 a2 = 0.42385546 rdsw = 65.968
+ rdswmin = 0 rdw = 0 rdwmin = 0
+ rsw = 0 rswmin = 0 prwb = 0
+ prwg = 0.021507 wr = 1 voff = -0.16985218591
+ wvoff = -3.603061541361336E-8 voffl = 5.8197729E-9 minv = 0
+ nfactor = 0.970603803870452 lnfactor = 3.128061320207972E-7 wnfactor = -6.126933424180614E-6
+ pnfactor = 7.026425502137226E-13 eta0 = 6.9413878E-4 etab = -0.054585923983
+ wetab = 1.01250411223112E-8 dsub = 0.45862506 cit = 0
+ cdsc = 0 cdscb = 0 cdscd = 9.344996332361596E-3
+ lcdscd = -9.19909385378762E-10 wcdscd = -6.974161118703411E-9 pcdscd = 8.796927868687733E-16
+ pclm = 0.910493994356733 lpclm = -9.291278866035492E-8 wpclm = -7.466974937914452E-7
+ ppclm = 8.885082736570152E-14 pdiblc1 = 0.35697215 pdiblc2 = 8.4061121E-3
+ pdiblcb = -0.10329577 drout = 0.50332666 pscbe1 = 7.9141988E8
+ pscbe2 = 1E-12 pvag = 0 delta = 0.01
+ fprout = 0 pdits = 0 pditsl = 0
+ pditsd = 0 lambda = 0 vtl = 0
+ lc = 5E-9 xn = 3 alpha0 = 5.090340648927998E-8
+ lalpha0 = -2.636672080931819E-15 walpha0 = -6.179636434294159E-14 palpha0 = 7.794746212761279E-21
+ alpha1 = 0.85 beta0 = 16.292709533605333 lbeta0 = -3.062491417990825E-7
+ wbeta0 = -1.191208802849842E-6 pbeta0 = 1.484713564335484E-13 aigbacc = 1
+ bigbacc = 0 cigbacc = 0 nigbacc = 0
+ aigbinv = 0.35 bigbinv = 0.03 cigbinv = 6E-3
+ eigbinv = 1.1 nigbinv = 0 aigc = 0.43
+ bigc = 0.054 cigc = 0.075 aigsd = 0.43
+ bigsd = 0.054 cigsd = 0.075 dlcig = 0
+ nigc = 0 poxedge = 1 pigcd = 1
+ ntox = 1 toxref = 4.148E-9 agidl = 0
+ bgidl = 2.3E9 cgidl = 0.5 egidl = 0.8
+ noia = 2.5E42 noib = 0 noic = 0
+ em = 4.1E7 af = 1 ef = 0.84
+ kf = 0 lintnoi = -1E-7 tnoia = 1.5E7
+ tnoib = 9.9E6 ntnoi = 1 rnoia = 0.94
+ rnoib = 0.26 xpart = 0 cgso = {2.449068E-10/sw_func_tox_lv_ratio}
+ cgdo = {2.449068E-10/sw_func_tox_lv_ratio} cgbo = {1E-13/sw_func_tox_lv_ratio} ckappas = 0.6
+ cf = 1.4067E-12 clc = 1E-7 cle = 0.6
+ dlc = 9.87908E-9 dwc = 0 vfbcv = -1
+ noff = 3.4037 voffcv = -0.17287 acde = 0.4
+ moin = 6.9 cgsl = {0/sw_func_tox_lv_ratio} cgdl = {0/sw_func_tox_lv_ratio}
+ ijthsrev = 0.1 ijthsfwd = 0.1 xjbvs = 1
+ bvs = 11.7 jss = 2.75E-3 jsws = 6E-10
+ cjs = {sw_nsd_pw_cj} mjs = 0.44 mjsws = 9E-4
+ cjsws = {3.67354204E-11*sw_func_nsd_pw_cj} cjswgs = {2.38232788E-10*sw_func_nsd_pw_cj} mjswgs = 0.8
+ pbs = 0.729 pbsws = 0.2 pbswgs = 0.95578
+ xrcrg1 = 12 xrcrg2 = 1 rbpb = 50
+ rbpd = 50 rbps = 50 rbdb = 50
+ rbsb = 50 gbmin = 1E-12 tnom = 30
+ ute = -1.3190432 kt1 = -0.215534954549333 lkt1 = -6.27779066888529E-9
+ wkt1 = -1.047286118636677E-7 pkt1 = 1.855891955419355E-14 kt1l = 0
+ kt2 = -0.028878939 ua1 = -2.3847336E-11 ub1 = 7.0775317E-19
+ uc1 = 1.4718625E-10 at = 1.359088031373332E5 lat = -8.277737580778665E-3
+ wat = 8.513157568891965E-3 pat = -4.639729888548389E-9 prt = 0
+ njs = 1.2928 xtis = 2 tpb = 1.2287E-3
+ tpbsw = 0 tpbswg = 0 tcj = 7.92E-4
+ tcjsw = 1E-5 tcjswg = 0 tvoff = 0
+ tvfbsdoff = 0 saref = 1.1E-6 sbref = 1.1E-6
+ wlod = 0 ku0 = -2.7E-8 kvsat = 0.2
+ kvth0 = 9.8E-9 tku0 = 0 llodku0 = 0
+ wlodku0 = 1 llodvth = 0 wlodvth = 1
+ lku0 = 0 wku0 = 0 pku0 = 0
+ lkvth0 = 0 wkvth0 = 2E-7 pkvth0 = 0
+ stk2 = 0 lodk2 = 1 steta0 = 0
+ lodeta0 = 1

.model nshort_model.33 nmos
+ level = 54 lmin = 8E-6 lmax = 2.02E-5 wmin = 5.5E-7
+ wmax = 1E-6 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 4.148E-9
+ toxm = 4.148E-9 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 9.999999999999999E22 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {2.1859E-8+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {1.1932E-8-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = 0 dwb = 0 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = 0.535717068985778 wvth0 = -8.23030700285759E-9
+ k1 = 0.442231847658844 wk1 = 2.99164526434649E-8 k2 = 0.017140093776693
+ wk2 = -1.559470917053764E-8 k3 = 2 k3b = 0.54
+ w0 = 0 lpe0 = 1.0325E-7 lpeb = -7.082E-8
+ vbm = -3 dvtp0 = 0 dvtp1 = 0
+ dvt0 = 0 dvt1 = 0.53 dvt2 = -0.032
+ dvt0w = -3.58 dvt1w = 1.6706E6 dvt2w = 0.068
+ vfbsdoff = 0 u0 = 0.029859968275111 wu0 = -1.222098058059803E-9
+ ua = -5.391390653933777E-10 wua = -1.1738111444639E-16 ub = 1.259250940445466E-18
+ wub = 1.035367090909283E-25 uc = 2.521508809333333E-11 wuc = 5.583844459310166E-19
+ ud = 0 up = 0 lp = 1
+ eu = 1.67 vsat = 8E4 a0 = 1.413124866231111
+ wa0 = -4.714744352521944E-8 ags = 0.304713571897778 wags = 3.86275082124493E-8
+ b0 = -2.472231259555556E-8 wb0 = 2.364150253350306E-14 b1 = -2.212902368444445E-9
+ wb1 = 2.116158702700791E-15 keta = 5.049480961619115E-3 wketa = -6.295050121010449E-9
+ a1 = 0 a2 = 0.42385546 rdsw = 65.968
+ rdswmin = 0 rdw = 0 rdwmin = 0
+ rsw = 0 rswmin = 0 prwb = 0
+ prwg = 0.021507 wr = 1 voff = -0.103792223045867
+ wvoff = -7.291790779592537E-9 voffl = 5.8197729E-9 minv = 0
+ nfactor = 2.985191588888889 wnfactor = -6.186340200584457E-8 eta0 = 0.08
+ etab = -0.07 dsub = 0.56 cit = 0
+ cdsc = 0 cdscb = 0 cdscd = 5.4E-3
+ pclm = 0.113520895537778 wpclm = -2.867879728465721E-8 pdiblc1 = 0.39
+ pdiblc2 = 4.922590564592E-3 wpdiblc2 = -1.694740043987767E-9 pdiblcb = -4.686452285863112
+ wpdiblcb = 2.360009386191348E-6 drout = 0.56 pscbe1 = 8.588488658986223E8
+ wpscbe1 = -93.07977148766628 pscbe2 = 1E-12 pvag = 0
+ delta = 0.01 fprout = 0 pdits = 0
+ pditsl = 0 pditsd = 0 lambda = 0
+ vtl = 0 lc = 5E-9 xn = 3
+ alpha0 = 3E-8 alpha1 = 0.85 beta0 = 13.86
+ aigbacc = 1 bigbacc = 0 cigbacc = 0
+ nigbacc = 0 aigbinv = 0.35 bigbinv = 0.03
+ cigbinv = 6E-3 eigbinv = 1.1 nigbinv = 0
+ aigc = 0.43 bigc = 0.054 cigc = 0.075
+ aigsd = 0.43 bigsd = 0.054 cigsd = 0.075
+ dlcig = 0 nigc = 0 poxedge = 1
+ pigcd = 1 ntox = 1 toxref = 4.148E-9
+ agidl = 0 bgidl = 2.3E9 cgidl = 0.5
+ egidl = 0.8 noia = 2.5E42 noib = 0
+ noic = 0 em = 4.1E7 af = 1
+ ef = 0.84 kf = 0 lintnoi = -1E-7
+ tnoia = 1.5E7 tnoib = 9.9E6 ntnoi = 1
+ rnoia = 0.94 rnoib = 0.26 xpart = 0
+ cgso = {2.449068E-10/sw_func_tox_lv_ratio} cgdo = {2.449068E-10/sw_func_tox_lv_ratio} cgbo = {1E-13/sw_func_tox_lv_ratio}
+ ckappas = 0.6 cf = 1.4067E-12 clc = 1E-7
+ cle = 0.6 dlc = 9.87908E-9 dwc = 0
+ vfbcv = -1 noff = 3.4037 voffcv = -0.17287
+ acde = 0.4 moin = 6.9 cgsl = {0/sw_func_tox_lv_ratio}
+ cgdl = {0/sw_func_tox_lv_ratio} ijthsrev = 0.1 ijthsfwd = 0.1
+ xjbvs = 1 bvs = 11.7 jss = 2.75E-3
+ jsws = 6E-10 cjs = {sw_nsd_pw_cj} mjs = 0.44
+ mjsws = 9E-4 cjsws = {3.67354204E-11*sw_func_nsd_pw_cj} cjswgs = {2.38232788E-10*sw_func_nsd_pw_cj}
+ mjswgs = 0.8 pbs = 0.729 pbsws = 0.2
+ pbswgs = 0.95578 xrcrg1 = 12 xrcrg2 = 1
+ rbpb = 50 rbpd = 50 rbps = 50
+ rbdb = 50 rbsb = 50 gbmin = 1E-12
+ tnom = 30 ute = -1.313126607111111 wute = 2.431500670142775E-8
+ kt1 = -0.293987595288889 wkt1 = 1.441686238049253E-9 kt1l = 0
+ kt2 = -0.020710160521044 wkt2 = 7.029296295742312E-11 ua1 = 1.461044291111111E-9
+ wua1 = -1.027470415923155E-16 ub1 = -1.045060260222222E-18 wub1 = 9.849729484582725E-26
+ uc1 = -2.984207669519112E-11 wuc1 = 5.196200851144749E-18 at = 1.4E5
+ prt = 0 njs = 1.2928 xtis = 2
+ tpb = 1.2287E-3 tpbsw = 0 tpbswg = 0
+ tcj = 7.92E-4 tcjsw = 1E-5 tcjswg = 0
+ tvoff = 0 tvfbsdoff = 0 saref = 3E-6
+ sbref = 3E-6 wlod = 0 ku0 = -2.7E-8
+ kvsat = 0.2 kvth0 = 9.8E-9 tku0 = 0
+ llodku0 = 0 wlodku0 = 1 llodvth = 0
+ wlodvth = 1 lku0 = 0 wku0 = 0
+ pku0 = 0 lkvth0 = 0 wkvth0 = 2E-7
+ pkvth0 = 0 stk2 = 0 lodk2 = 1
+ steta0 = 0 lodeta0 = 1

.model nshort_model.34 nmos
+ level = 54 lmin = 4E-6 lmax = 8E-6 wmin = 5.5E-7
+ wmax = 1E-6 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 4.148E-9
+ toxm = 4.148E-9 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 9.999999999999999E22 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {2.1859E-8+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {1.1932E-8-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = 0 dwb = 0 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = 0.533989010007646 lvth0 = 1.378323342560346E-8
+ wvth0 = -1.115615351062776E-8 pvth0 = 2.333694966109995E-14 k1 = 0.4793017487653
+ lk1 = -2.956745727316402E-7 wk1 = -2.144285892777418E-8 pk1 = 4.096488539585766E-13
+ k2 = 3.211561506779391E-3 lk2 = 1.110958676652188E-7 wk2 = 5.861465150105437E-9
+ pk2 = -1.711373644211568E-13 k3 = 2 k3b = 0.54
+ w0 = 0 lpe0 = 1.0325E-7 lpeb = -7.082E-8
+ vbm = -3 dvtp0 = 0 dvtp1 = 0
+ dvt0 = 0 dvt1 = 0.53 dvt2 = -0.032
+ dvt0w = -3.58 dvt1w = 1.6706E6 dvt2w = 0.068
+ vfbsdoff = 0 u0 = 0.033207448184829 lu0 = -2.669995501717692E-8
+ wu0 = -3.791384427775018E-9 pu0 = 2.049297750779484E-14 ua = -2.286659081973656E-10
+ lua = -2.476376126144771E-15 wua = -3.787969334888164E-16 pua = 2.085088125233783E-21
+ ub = 1.059282761648736E-18 lub = 1.594973389755044E-24 wub = 2.878881074732996E-25
+ pub = -1.470411825287973E-30 uc = 4.49161968717749E-11 luc = -1.571387229676438E-16
+ wuc = -1.788028784022451E-17 puc = 1.470693578138074E-22 ud = 0
+ up = 0 lp = 1 eu = 1.67
+ vsat = 8E4 a0 = 1.585871130159841 la0 = -1.377847694587445E-6
+ wa0 = -8.931223057666468E-8 pa0 = 3.363120759333663E-13 ags = 0.345633281829748
+ lags = -3.263811714979435E-7 wags = 7.764843353457575E-9 pags = 2.461648122377388E-13
+ b0 = -1.217879875970887E-8 lb0 = -1.000487722725949E-13 wb0 = 1.164636603553192E-14
+ pb0 = 9.567484004638159E-20 b1 = -6.731457841725369E-10 lb1 = -1.22813079230482E-14
+ wb1 = 6.437171967800818E-16 pb1 = 1.174439370326838E-20 keta = -7.466520972306588E-3
+ lketa = 9.98293336012544E-8 wketa = -5.061495458800998E-9 pketa = -9.838999749216645E-15
+ a1 = 0 a2 = 0.42385546 rdsw = 65.968
+ rdswmin = 0 rdw = 0 rdwmin = 0
+ rsw = 0 rswmin = 0 prwb = 0
+ prwg = 0.021507 wr = 1 voff = -0.115435468609223
+ lvoff = 9.286811009472848E-8 wvoff = -1.297495098160795E-9 pvoff = -4.781131757931225E-14
+ voffl = 5.8197729E-9 minv = 0 nfactor = 3.077439013950453
+ lnfactor = -7.357780079408492E-7 wnfactor = -1.22416168630357E-7 pnfactor = 4.829771017733717E-13
+ eta0 = 0.08 etab = -0.07 dsub = 0.56
+ cit = 0 cdsc = 0 cdscb = 0
+ cdscd = 5.4E-3 pclm = 9.145618255666621E-3 lpclm = 8.325114066398302E-7
+ wpclm = -3.562735040885561E-7 ppclm = 2.612939934348023E-12 pdiblc1 = 0.39
+ pdiblc2 = 8.133287302480884E-3 lpdiblc2 = -2.56089538361581E-8 wpdiblc2 = -4.949739150442705E-9
+ ppdiblc2 = 2.596231555296306E-14 pdiblcb = -9.320094347388764 lpdiblcb = 3.695855925804898E-5
+ wpdiblcb = 4.705938956384679E-6 ppdiblcb = -1.871145329828355E-11 drout = 0.56
+ pscbe1 = 9.33738594770141E8 lpscbe1 = -597.3306624823596 wpscbe1 = -149.21504247977285
+ ppscbe1 = 4.477425558298969E-4 pscbe2 = 1E-12 pvag = 0
+ delta = 0.01 fprout = 0 pdits = 0
+ pditsl = 0 pditsd = 0 lambda = 0
+ vtl = 0 lc = 5E-9 xn = 3
+ alpha0 = 3E-8 alpha1 = 0.85 beta0 = 13.86
+ aigbacc = 1 bigbacc = 0 cigbacc = 0
+ nigbacc = 0 aigbinv = 0.35 bigbinv = 0.03
+ cigbinv = 6E-3 eigbinv = 1.1 nigbinv = 0
+ aigc = 0.43 bigc = 0.054 cigc = 0.075
+ aigsd = 0.43 bigsd = 0.054 cigsd = 0.075
+ dlcig = 0 nigc = 0 poxedge = 1
+ pigcd = 1 ntox = 1 toxref = 4.148E-9
+ agidl = 0 bgidl = 2.3E9 cgidl = 0.5
+ egidl = 0.8 noia = 2.5E42 noib = 0
+ noic = 0 em = 4.1E7 af = 1
+ ef = 0.84 kf = 0 lintnoi = -1E-7
+ tnoia = 1.5E7 tnoib = 9.9E6 ntnoi = 1
+ rnoia = 0.94 rnoib = 0.26 xpart = 0
+ cgso = {2.449068E-10/sw_func_tox_lv_ratio} cgdo = {2.449068E-10/sw_func_tox_lv_ratio} cgbo = {1E-13/sw_func_tox_lv_ratio}
+ ckappas = 0.6 cf = 1.4067E-12 clc = 1E-7
+ cle = 0.6 dlc = 9.87908E-9 dwc = 0
+ vfbcv = -1 noff = 3.4037 voffcv = -0.17287
+ acde = 0.4 moin = 6.9 cgsl = {0/sw_func_tox_lv_ratio}
+ cgdl = {0/sw_func_tox_lv_ratio} ijthsrev = 0.1 ijthsfwd = 0.1
+ xjbvs = 1 bvs = 11.7 jss = 2.75E-3
+ jsws = 6E-10 cjs = {sw_nsd_pw_cj} mjs = 0.44
+ mjsws = 9E-4 cjsws = {3.67354204E-11*sw_func_nsd_pw_cj} cjswgs = {2.38232788E-10*sw_func_nsd_pw_cj}
+ mjswgs = 0.8 pbs = 0.729 pbsws = 0.2
+ pbswgs = 0.95578 xrcrg1 = 12 xrcrg2 = 1
+ rbpb = 50 rbpd = 50 rbps = 50
+ rbdb = 50 rbsb = 50 gbmin = 1E-12
+ tnom = 30 ute = -1.778612170479028 lute = 3.712776159459118E-6
+ wute = 2.772438388849316E-7 pute = -2.017394763816804E-12 kt1 = -0.296869310767173
+ lkt1 = 2.298495456810108E-8 wkt1 = 5.366628369607223E-9 pkt1 = -3.130587223343625E-14
+ kt1l = 0 kt2 = -0.032703727713221 lkt2 = 9.56623230499375E-8
+ wkt2 = 1.1598198788362E-8 pkt2 = -9.194814465861916E-14 ua1 = 9.55745060569633E-10
+ lua1 = 4.030335383494182E-15 wua1 = 2.835977390685328E-16 pua1 = -3.081538513441097E-21
+ ub1 = -8.328632257334639E-19 lub1 = -1.692512405879028E-24 wub1 = -9.851982762709029E-26
+ pub1 = 1.571435363172647E-30 uc1 = 1.530361460488377E-11 luc1 = -3.600881736234139E-16
+ wuc1 = -4.379667969058942E-17 puc1 = 3.907738782326254E-22 at = 1.4E5
+ prt = 0 njs = 1.2928 xtis = 2
+ tpb = 1.2287E-3 tpbsw = 0 tpbswg = 0
+ tcj = 7.92E-4 tcjsw = 1E-5 tcjswg = 0
+ tvoff = 0 tvfbsdoff = 0 saref = 3E-6
+ sbref = 3E-6 wlod = 0 ku0 = -2.7E-8
+ kvsat = 0.2 kvth0 = 9.8E-9 tku0 = 0
+ llodku0 = 0 wlodku0 = 1 llodvth = 0
+ wlodvth = 1 lku0 = 0 wku0 = 0
+ pku0 = 0 lkvth0 = 0 wkvth0 = 2E-7
+ pkvth0 = 0 stk2 = 0 lodk2 = 1
+ steta0 = 0 lodeta0 = 1

.model nshort_model.35 nmos
+ level = 54 lmin = 2E-6 lmax = 4E-6 wmin = 5.5E-7
+ wmax = 1E-6 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 4.148E-9
+ toxm = 4.148E-9 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 9.999999999999999E22 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {2.1859E-8+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {1.1932E-8-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = 0 dwb = 0 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = 0.479816508865313 lvth0 = 2.291804654276729E-7
+ wvth0 = 2.826373854344638E-8 pvth0 = -1.334019022512182E-13 k1 = 0.309497854226312
+ lk1 = 3.794888052850331E-7 wk1 = 1.263947088694731E-7 pk1 = -1.781734215124992E-13
+ k2 = 0.080082763758251 lk2 = -1.945544869701378E-7 wk2 = -6.064703668853995E-8
+ pk2 = 9.33094840455474E-14 k3 = 2 k3b = 0.54
+ w0 = 0 lpe0 = 1.0325E-7 lpeb = -7.082E-8
+ vbm = -3 dvtp0 = 0 dvtp1 = 0
+ dvt0 = 0 dvt1 = 0.53 dvt2 = -0.032
+ dvt0w = -3.58 dvt1w = 1.6706E6 dvt2w = 0.068
+ vfbsdoff = 0 u0 = 0.028279900951863 lu0 = -7.10735707248039E-9
+ wu0 = 9.205508792440144E-10 pu0 = 1.757681903885414E-15 ua = 2.680915076921181E-10
+ lua = -4.451551170729919E-15 wua = -4.929216170526986E-16 pua = 2.538863388040743E-21
+ ub = -1.365293846439406E-19 lub = 6.349685113866622E-24 wub = 9.170270030734071E-25
+ pub = -3.971953637083803E-30 uc = -4.639433909702059E-11 luc = 2.059243862771788E-16
+ wuc = 4.149976071729185E-17 puc = -8.903379093748147E-23 ud = 0
+ up = 0 lp = 1 eu = 1.67
+ vsat = 8E4 a0 = 1.222055957833506 la0 = 6.873090944550226E-8
+ wa0 = 1.967147753875323E-7 pa0 = -8.00970199453092E-13 ags = 8.706105517577833E-3
+ lags = 1.013287103615222E-6 wags = 1.610392596960605E-7 pags = -3.632751124610728E-13
+ b0 = -7.256891108198214E-10 lb0 = -1.4558789385949E-13 wb0 = 6.939634342729998E-16
+ pb0 = 1.392230823157408E-19 b1 = 1.469731719988644E-9 lb1 = -2.080168031093363E-14
+ wb1 = -1.405477988654182E-15 pb1 = 1.989227245110023E-20 keta = 0.059219497364668
+ lketa = -1.653233446050501E-7 wketa = -2.97195507760595E-8 pketa = 8.820478168772631E-14
+ a1 = 0 a2 = 0.42385546 rdsw = 65.968
+ rdswmin = 0 rdw = 0 rdwmin = 0
+ rsw = 0 rswmin = 0 prwb = 0
+ prwg = 0.021507 wr = 1 voff = -0.029221150718578
+ lvoff = -2.49931742985711E-7 wvoff = -5.468761251889512E-8 pvoff = 1.644750503414966E-13
+ voffl = 5.8197729E-9 minv = 0 nfactor = 4.333058725516963
+ lnfactor = -5.72829274541006E-6 wnfactor = -9.073070698962012E-7 pnfactor = 3.60381007036894E-12
+ eta0 = -8.375917627759966E-3 leta0 = 3.513946676127711E-7 weta0 = 8.451229926090958E-8
+ peta0 = -3.36032395534076E-13 etab = 7.259450001626699E-3 letab = -3.07194080491668E-7
+ wetab = -7.388182136645556E-8 petab = 2.937641696807332E-13 dsub = 0.226505971216
+ ldsub = 1.326017613633099E-6 wdsub = 3.189143368336211E-7 pdsub = -1.268046775600287E-12
+ cit = 0 cdsc = 0 cdscb = 0
+ cdscd = 5.4E-3 pclm = -0.173199213742234 lpclm = 1.557539257560636E-6
+ wpclm = 6.528678232146496E-7 ppclm = -1.399543226230037E-12 pdiblc1 = 0.39
+ pdiblc2 = 2.247446357645484E-4 lpdiblc2 = 5.836487368508731E-9 wpdiblc2 = 1.138852495148438E-9
+ ppdiblc2 = 1.753247121628876E-15 pdiblcb = -0.011104415467333 lpdiblcb = -5.525073390137912E-8
+ wpdiblcb = -1.328809736806755E-8 ppdiblcb = 5.283528231667863E-14 drout = 0.56
+ pscbe1 = 7.672160893863049E8 lpscbe1 = 64.78546598450512 wpscbe1 = -72.77837315772861
+ ppscbe1 = 1.438199632184212E-4 pscbe2 = 1E-12 pvag = 0
+ delta = 0.01 fprout = 0 pdits = 0
+ pditsl = 0 pditsd = 0 lambda = 0
+ vtl = 0 lc = 5E-9 xn = 3
+ alpha0 = 3E-8 alpha1 = 0.85 beta0 = 13.86
+ aigbacc = 1 bigbacc = 0 cigbacc = 0
+ nigbacc = 0 aigbinv = 0.35 bigbinv = 0.03
+ cigbinv = 6E-3 eigbinv = 1.1 nigbinv = 0
+ aigc = 0.43 bigc = 0.054 cigc = 0.075
+ aigsd = 0.43 bigsd = 0.054 cigsd = 0.075
+ dlcig = 0 nigc = 0 poxedge = 1
+ pigcd = 1 ntox = 1 toxref = 4.148E-9
+ agidl = 0 bgidl = 2.3E9 cgidl = 0.5
+ egidl = 0.8 noia = 2.5E42 noib = 0
+ noic = 0 em = 4.1E7 af = 1
+ ef = 0.84 kf = 0 lintnoi = -1E-7
+ tnoia = 1.5E7 tnoib = 9.9E6 ntnoi = 1
+ rnoia = 0.94 rnoib = 0.26 xpart = 0
+ cgso = {2.449068E-10/sw_func_tox_lv_ratio} cgdo = {2.449068E-10/sw_func_tox_lv_ratio} cgbo = {1E-13/sw_func_tox_lv_ratio}
+ ckappas = 0.6 cf = 1.4067E-12 clc = 1E-7
+ cle = 0.6 dlc = 9.87908E-9 dwc = 0
+ vfbcv = -1 noff = 3.4037 voffcv = -0.17287
+ acde = 0.4 moin = 6.9 cgsl = {0/sw_func_tox_lv_ratio}
+ cgdl = {0/sw_func_tox_lv_ratio} ijthsrev = 0.1 ijthsfwd = 0.1
+ xjbvs = 1 bvs = 11.7 jss = 2.75E-3
+ jsws = 6E-10 cjs = {sw_nsd_pw_cj} mjs = 0.44
+ mjsws = 9E-4 cjsws = {3.67354204E-11*sw_func_nsd_pw_cj} cjswgs = {2.38232788E-10*sw_func_nsd_pw_cj}
+ mjswgs = 0.8 pbs = 0.729 pbsws = 0.2
+ pbswgs = 0.95578 xrcrg1 = 12 xrcrg2 = 1
+ rbpb = 50 rbpd = 50 rbps = 50
+ rbdb = 50 rbsb = 50 gbmin = 1E-12
+ tnom = 30 ute = -2.716140923075198 lute = 7.44051798369184E-6
+ wute = 9.328743176252128E-7 pute = -4.62427071303327E-12 kt1 = -0.337349019970748
+ lkt1 = 1.839377836019658E-7 wkt1 = 3.981311986001949E-8 pkt1 = -1.682698071221581E-13
+ kt1l = 0 kt2 = -0.033676888860133 lkt2 = 9.953174411997703E-8
+ wkt2 = 9.576883120965799E-9 pkt2 = -8.39111186661211E-14 ua1 = -3.840292346504822E-9
+ lua1 = 2.310003237510958E-14 wua1 = 3.02788353132741E-15 pua1 = -1.399319204633014E-20
+ ub1 = 3.410975448946843E-18 lub1 = -1.856659213846768E-23 wub1 = -2.479303599426119E-24
+ pub1 = 1.103775542643855E-29 uc1 = -2.326720172007665E-11 luc1 = -2.067253622843512E-16
+ wuc1 = 1.604126213163065E-17 puc1 = 1.528500835873906E-22 at = 1.664220448244176E5
+ lat = -0.10505764361998 wat = 1.945377454685089E-3 pat = -7.73508533116175E-9
+ prt = 0 njs = 1.2928 xtis = 2
+ tpb = 1.2287E-3 tpbsw = 0 tpbswg = 0
+ tcj = 7.92E-4 tcjsw = 1E-5 tcjswg = 0
+ tvoff = 0 tvfbsdoff = 0 saref = 3E-6
+ sbref = 3E-6 wlod = 0 ku0 = -2.7E-8
+ kvsat = 0.2 kvth0 = 9.8E-9 tku0 = 0
+ llodku0 = 0 wlodku0 = 1 llodvth = 0
+ wlodvth = 1 lku0 = 0 wku0 = 0
+ pku0 = 0 lkvth0 = 0 wkvth0 = 2E-7
+ pkvth0 = 0 stk2 = 0 lodk2 = 1
+ steta0 = 0 lodeta0 = 1

.model nshort_model.36 nmos
+ level = 54 lmin = 1E-6 lmax = 2E-6 wmin = 5.5E-7
+ wmax = 1E-6 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 4.148E-9
+ toxm = 4.148E-9 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 9.999999999999999E22 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {2.1859E-8+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {1.1932E-8-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = 0 dwb = 0 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = 0.57447160566449 lvth0 = 4.212912105933517E-8
+ wvth0 = -4.543095872824798E-8 pvth0 = 1.222884203647877E-14 k1 = 0.60554879394503
+ lk1 = -2.055481145269547E-7 wk1 = -7.083494066279599E-9 pk1 = 8.559766052414735E-14
+ k2 = -0.050893092144031 lk2 = 6.427161700917363E-8 wk2 = 4.524174599334751E-10
+ pk2 = -2.743134687760028E-14 k3 = 2 k3b = 0.54
+ w0 = 0 lpe0 = 1.0325E-7 lpeb = -7.082E-8
+ vbm = -3 dvtp0 = 0 dvtp1 = 0
+ dvt0 = 0 dvt1 = 0.53 dvt2 = -0.032
+ dvt0w = -3.58 dvt1w = 1.6706E6 dvt2w = 0.068
+ vfbsdoff = 0 u0 = 0.026057446902643 lu0 = -2.715485617470194E-9
+ wu0 = 2.429468205836287E-9 pu0 = -1.224143946217334E-15 ua = -2.281103302137393E-9
+ lua = 5.860044639873304E-16 wua = 1.294334143309266E-15 pua = -9.929970612179069E-22
+ ub = 3.71385621772816E-18 lub = -1.259200488862569E-24 wub = -1.849135549566848E-24
+ pub = 1.494359765040499E-30 uc = 1.217705713713993E-11 luc = 9.017934160858975E-17
+ wuc = 2.510236430883195E-17 puc = -5.663030558845315E-23 ud = 0
+ up = 0 lp = 1 eu = 1.67
+ vsat = 6.300794362546317E4 lvsat = 0.033578614315752 wvsat = 6.914584790434821E-3
+ pvsat = -1.36641599294307E-8 a0 = 2.448401097977582 la0 = -2.354693870418253E-6
+ wa0 = -9.87414241758517E-7 pa0 = 1.539029779973833E-12 ags = 1.008765531036257
+ lags = -9.629663292915569E-7 wags = -6.517902484816878E-7 pags = 1.24298654051127E-12
+ b0 = -2.162691899247486E-8 lb0 = -1.042842210460757E-13 wb0 = 2.068143334796185E-14
+ pb0 = 9.972512347038337E-20 b1 = -1.547768692594276E-8 lb1 = 1.268872378236267E-14
+ wb1 = 1.480103340891439E-14 pb1 = -1.213399815604534E-20 keta = -0.136920506745836
+ lketa = 2.222759785578639E-7 wketa = 1.053185851803794E-7 pketa = -1.786489401486871E-13
+ a1 = 0 a2 = 0.42385546 rdsw = 65.968
+ rdswmin = 0 rdw = 0 rdwmin = 0
+ rsw = 0 rswmin = 0 prwb = 0
+ prwg = 0.021507 wr = 1 voff = -0.14163685757588
+ lvoff = -2.778301769954952E-8 wvoff = 3.88939985659726E-8 pvoff = -2.045494026130949E-14
+ voffl = 5.8197729E-9 minv = 0 nfactor = 1.938035751111073
+ lnfactor = -9.954016248595036E-7 wnfactor = 8.410181577716368E-7 pnfactor = 1.488816482663299E-13
+ eta0 = 0.332371767287599 leta0 = -3.219690994651274E-7 weta0 = -1.690245460113029E-7
+ peta0 = 1.649908917347728E-13 etab = -0.210486945003253 letab = 1.231024095476958E-7
+ wetab = 1.477636427329112E-7 petab = -1.44237411162733E-13 dsub = 1.519828857568001
+ ldsub = -1.229764301710998E-6 wdsub = -6.378286736672425E-7 pdsub = 6.226075301988474E-13
+ cit = 0 cdsc = 0 cdscb = 0
+ cdscd = 5.4E-3 pclm = 0.743299311994367 lpclm = -2.535864730943879E-7
+ wpclm = -3.005574032877065E-7 ppclm = 4.84554687169423E-13 pdiblc1 = 0.457273537408558
+ lpdiblc1 = -1.329416591203989E-7 wpdiblc1 = -1.645022150141637E-8 ppdiblc1 = 3.250787491692294E-14
+ pdiblc2 = -6.087635397317775E-4 lpdiblc2 = 7.483612880401338E-9 wpdiblc2 = 5.171651582822114E-9
+ ppdiblc2 = -6.216112336290233E-15 pdiblcb = 0.025011463129838 lpdiblcb = -1.266206217688786E-7
+ wpdiblcb = -2.5074239444662E-8 ppdiblcb = 7.612630197535167E-14 drout = 1.292532976204963
+ ldrout = -1.447584785465771E-6 wdrout = -5.486337709041196E-7 pdrout = 1.084174945499383E-12
+ pscbe1 = 7.274043684930816E8 lpscbe1 = 143.45884086355582 wpscbe1 = 69.42189568869902
+ ppscbe1 = -1.371871072586829E-4 pscbe2 = 1E-12 pvag = 0
+ delta = 0.01 fprout = 0 pdits = 0
+ pditsl = 0 pditsd = 0 lambda = 0
+ vtl = 0 lc = 5E-9 xn = 3
+ alpha0 = 6.061730283591342E-6 lalpha0 = -1.191951935569506E-11 walpha0 = -5.766914945509673E-12
+ palpha0 = 1.13962082327597E-17 alpha1 = 1.16737683735968 lalpha1 = -6.271797938726093E-7
+ walpha1 = -1.606821799721337E-7 palpha1 = 3.175298404014124E-13 beta0 = 17.817993580472464
+ lbeta0 = -7.821533602140531E-6 wbeta0 = -3.784958017121369E-6 pbeta0 = 7.479591796122151E-12
+ aigbacc = 1 bigbacc = 0 cigbacc = 0
+ nigbacc = 0 aigbinv = 0.35 bigbinv = 0.03
+ cigbinv = 6E-3 eigbinv = 1.1 nigbinv = 0
+ aigc = 0.43 bigc = 0.054 cigc = 0.075
+ aigsd = 0.43 bigsd = 0.054 cigsd = 0.075
+ dlcig = 0 nigc = 0 poxedge = 1
+ pigcd = 1 ntox = 1 toxref = 4.148E-9
+ agidl = 0 bgidl = 2.3E9 cgidl = 0.5
+ egidl = 0.8 noia = 2.5E42 noib = 0
+ noic = 0 em = 4.1E7 af = 1
+ ef = 0.84 kf = 0 lintnoi = -1E-7
+ tnoia = 1.5E7 tnoib = 9.9E6 ntnoi = 1
+ rnoia = 0.94 rnoib = 0.26 xpart = 0
+ cgso = {2.449068E-10/sw_func_tox_lv_ratio} cgdo = {2.449068E-10/sw_func_tox_lv_ratio} cgbo = {1E-13/sw_func_tox_lv_ratio}
+ ckappas = 0.6 cf = 1.4067E-12 clc = 1E-7
+ cle = 0.6 dlc = 9.87908E-9 dwc = 0
+ vfbcv = -1 noff = 3.4037 voffcv = -0.17287
+ acde = 0.4 moin = 6.9 cgsl = {0/sw_func_tox_lv_ratio}
+ cgdl = {0/sw_func_tox_lv_ratio} ijthsrev = 0.1 ijthsfwd = 0.1
+ xjbvs = 1 bvs = 11.7 jss = 2.75E-3
+ jsws = 6E-10 cjs = {sw_nsd_pw_cj} mjs = 0.44
+ mjsws = 9E-4 cjsws = {3.67354204E-11*sw_func_nsd_pw_cj} cjswgs = {2.38232788E-10*sw_func_nsd_pw_cj}
+ mjswgs = 0.8 pbs = 0.729 pbsws = 0.2
+ pbswgs = 0.95578 xrcrg1 = 12 xrcrg2 = 1
+ rbpb = 50 rbpd = 50 rbps = 50
+ rbdb = 50 rbsb = 50 gbmin = 1E-12
+ tnom = 30 ute = 3.064332053459886 lute = -3.982482762266291E-6
+ wute = -2.751578156378582E-6 pute = 2.656708461134692E-12 kt1 = -0.251980911486516
+ lkt1 = 1.52387911743705E-8 wkt1 = -7.067200723562515E-8 pkt1 = 5.006382999612067E-14
+ kt1l = 0 kt2 = 0.078338823843009 lkt2 = -1.2182653831836E-7
+ wkt2 = -7.454382573878319E-8 pkt2 = 8.232284245714783E-14 ua1 = 1.433326139777934E-8
+ lua1 = -1.281338142690514E-14 wua1 = -8.046716593140549E-15 pua1 = 7.891723945235472E-21
+ ub1 = -1.096972014418296E-17 lub1 = 9.851618128157481E-24 wub1 = 6.036067237561389E-24
+ pub1 = -5.789775437882594E-30 uc1 = -2.450958859913201E-10 luc1 = 2.316382865366869E-16
+ wuc1 = 1.604278017359051E-16 puc1 = -1.324773552400419E-22 at = 1.148567185279983E5
+ lat = -3.15754597387968E-3 wat = 0.020292406775289 pat = -4.399131046466354E-8
+ prt = 0 njs = 1.2928 xtis = 2
+ tpb = 1.2287E-3 tpbsw = 0 tpbswg = 0
+ tcj = 7.92E-4 tcjsw = 1E-5 tcjswg = 0
+ tvoff = 0 tvfbsdoff = 0 saref = 3E-6
+ sbref = 3E-6 wlod = 0 ku0 = -2.7E-8
+ kvsat = 0.2 kvth0 = 9.8E-9 tku0 = 0
+ llodku0 = 0 wlodku0 = 1 llodvth = 0
+ wlodvth = 1 lku0 = 0 wku0 = 0
+ pku0 = 0 lkvth0 = 0 wkvth0 = 2E-7
+ pkvth0 = 0 stk2 = 0 lodk2 = 1
+ steta0 = 0 lodeta0 = 1

.model nshort_model.37 nmos
+ level = 54 lmin = 5E-7 lmax = 1E-6 wmin = 5.5E-7
+ wmax = 1E-6 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 4.148E-9
+ toxm = 4.148E-9 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 9.999999999999999E22 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {2.1859E-8+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {1.1932E-8-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = 0 dwb = 0 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = 0.642181684593901 lvth0 = -2.396512454650492E-8
+ wvth0 = -5.276382311347358E-8 pvth0 = 1.938671494601536E-14 k1 = 0.139684346858981
+ lk1 = 2.491989433938325E-7 wk1 = 2.480422126526219E-7 pk1 = -1.634397263296143E-13
+ k2 = 0.090863259697772 lk2 = -7.410186125227674E-8 wk2 = -8.06074465417255E-8
+ pk2 = 5.169410452952311E-14 k3 = 2 k3b = 0.54
+ w0 = 0 lpe0 = 1.0325E-7 lpeb = -7.082E-8
+ vbm = -3 dvtp0 = 0 dvtp1 = 0
+ dvt0 = 0 dvt1 = 0.53 dvt2 = -0.032
+ dvt0w = -3.58 dvt1w = 1.6706E6 dvt2w = 0.068
+ vfbsdoff = 0 u0 = 0.023807246563211 lu0 = -5.18984058938396E-10
+ wu0 = 2.911977439785111E-9 pu0 = -1.695138579807203E-15 ua = -1.830461650157239E-9
+ lua = 1.461169243900316E-16 wua = 5.062942961165194E-16 pua = -2.237629969385683E-22
+ ub = 2.793480054008978E-18 lub = -3.607881819143823E-25 wub = -5.541379369174536E-25
+ pub = 2.302659754193703E-31 uc = 1.035048829792666E-10 luc = 1.030963002359616E-18
+ wuc = -3.863750957289777E-17 puc = 5.588479942962971E-24 ud = 0
+ up = 0 lp = 1 eu = 1.67
+ vsat = 1.222114358694848E5 lvsat = -0.024212045789359 wvsat = -0.06231274609256
+ pvsat = 5.391112992937248E-8 a0 = -1.481487359441263 la0 = 1.481411728852749E-6
+ wa0 = 1.268589768631483E-6 pa0 = -6.631369507122203E-13 ags = -2.005442603865723
+ lags = 1.979310742679121E-6 wags = 2.175488743765346E-6 pags = -1.516822265864781E-12
+ b0 = -2.507900704874283E-7 lb0 = 1.194101810016022E-13 wb0 = 2.398260301858589E-13
+ pb0 = -1.141898067085741E-19 b1 = -4.839207245558785E-9 lb1 = 2.304120781071377E-15
+ wb1 = 4.627646783197446E-15 pb1 = -2.203389228764499E-21 keta = 0.233661609738782
+ lketa = -1.394625662989651E-7 wketa = -1.768201635200694E-7 pketa = 9.675684945277429E-14
+ a1 = 0 a2 = 0.42385546 rdsw = 65.968
+ rdswmin = 0 rdw = 0 rdwmin = 0
+ rsw = 0 rswmin = 0 prwb = 0
+ prwg = 0.021507 wr = 1 voff = -0.191649272984349
+ lvoff = 2.10359014276115E-8 wvoff = 3.31741162129793E-8 pvoff = -1.487155718078803E-14
+ voffl = 5.8197729E-9 minv = 0 nfactor = -1.338347778573884
+ lnfactor = 2.202794288273052E-6 wnfactor = 2.086603999591472E-6 pnfactor = -1.066979533024317E-12
+ eta0 = -0.461671384064159 leta0 = 4.531250061227721E-7 peta0 = 5.00042944074647E-20
+ etab = -0.1647601692866 letab = 7.846685760674456E-8 wetab = 3.201673127984144E-10
+ petab = -3.12526840045793E-16 dsub = 0.20592405551017 ldsub = 5.278547615052472E-8
+ wdsub = 3.123695738617558E-9 pdsub = -3.049151863511189E-15 cit = 0
+ cdsc = 0 cdscb = 0 cdscd = 5.4E-3
+ pclm = 0.416183988809078 lpclm = 6.572257001840719E-8 wpclm = 4.317119324795676E-7
+ ppclm = -2.302397731691008E-13 pdiblc1 = 0.374629793178768 lpdiblc1 = -5.227012520290875E-8
+ wpdiblc1 = 1.446641995924032E-7 ppdiblc1 = -1.247617116319137E-13 pdiblc2 = 0.010578902969153
+ lpdiblc2 = -3.437071154915309E-9 wpdiblc2 = -7.381156845624805E-10 ppdiblc2 = -4.473757549745034E-16
+ pdiblcb = -0.25517845695896 lpdiblcb = 1.468828460669207E-7 wpdiblcb = 1.746138700974975E-7
+ ppdiblcb = -1.187964505206937E-13 drout = -1.324065739547297 ldrout = 1.106571418533777E-6
+ wdrout = 1.097267644261779E-6 pdrout = -5.224486782949962E-13 pscbe1 = 5.562258316060067E8
+ lpscbe1 = 310.55237314635747 wpscbe1 = 233.11684930014468 ppscbe1 = -2.96975644497145E-4
+ pscbe2 = 1E-12 pvag = 0 delta = 0.01
+ fprout = 0 pdits = 0 pditsl = 0
+ pditsd = 0 lambda = 0 vtl = 0
+ lc = 5E-9 xn = 3 alpha0 = -7.887244281928279E-6
+ lalpha0 = 1.696576880793002E-12 walpha0 = 7.568877889323694E-12 palpha0 = -1.621339241863201E-18
+ alpha1 = 0.21524632528064 lalpha1 = 3.022290756661772E-7 walpha1 = 3.213643599442671E-7
+ palpha1 = -1.530131408864236E-13 beta0 = 10.398784754840037 lbeta0 = -5.793767759229972E-7
+ wbeta0 = 3.309897837072059E-6 pbeta0 = 5.540475820331957E-13 aigbacc = 1
+ bigbacc = 0 cigbacc = 0 nigbacc = 0
+ aigbinv = 0.35 bigbinv = 0.03 cigbinv = 6E-3
+ eigbinv = 1.1 nigbinv = 0 aigc = 0.43
+ bigc = 0.054 cigc = 0.075 aigsd = 0.43
+ bigsd = 0.054 cigsd = 0.075 dlcig = 0
+ nigc = 0 poxedge = 1 pigcd = 1
+ ntox = 1 toxref = 4.148E-9 agidl = 0
+ bgidl = 2.3E9 cgidl = 0.5 egidl = 0.8
+ noia = 2.5E42 noib = 0 noic = 0
+ em = 4.1E7 af = 1 ef = 0.84
+ kf = 0 lintnoi = -1E-7 tnoia = 1.5E7
+ tnoib = 9.9E6 ntnoi = 1 rnoia = 0.94
+ rnoib = 0.26 xpart = 0 cgso = {2.449068E-10/sw_func_tox_lv_ratio}
+ cgdo = {2.449068E-10/sw_func_tox_lv_ratio} cgbo = {1E-13/sw_func_tox_lv_ratio} ckappas = 0.6
+ cf = 1.4067E-12 clc = 1E-7 cle = 0.6
+ dlc = 9.87908E-9 dwc = 0 vfbcv = -1
+ noff = 3.4037 voffcv = -0.17287 acde = 0.4
+ moin = 6.9 cgsl = {0/sw_func_tox_lv_ratio} cgdl = {0/sw_func_tox_lv_ratio}
+ ijthsrev = 0.1 ijthsfwd = 0.1 xjbvs = 1
+ bvs = 11.7 jss = 2.75E-3 jsws = 6E-10
+ cjs = {sw_nsd_pw_cj} mjs = 0.44 mjsws = 9E-4
+ cjsws = {3.67354204E-11*sw_func_nsd_pw_cj} cjswgs = {2.38232788E-10*sw_func_nsd_pw_cj} mjswgs = 0.8
+ pbs = 0.729 pbsws = 0.2 pbswgs = 0.95578
+ xrcrg1 = 12 xrcrg2 = 1 rbpb = 50
+ rbpd = 50 rbps = 50 rbdb = 50
+ rbsb = 50 gbmin = 1E-12 tnom = 30
+ ute = -0.905475277648852 lute = -1.074109133071304E-7 wute = 2.799069044982988E-8
+ pute = -5.652875473300725E-14 kt1 = -0.212389590849279 lkt1 = -2.340772218717955E-8
+ wkt1 = -2.945535738186284E-8 pkt1 = 9.830774274468547E-15 kt1l = 0
+ kt2 = -0.056493746119633 lkt2 = 9.788387194694128E-9 wkt2 = 1.949327233084588E-8
+ pkt2 = -9.470154304147621E-15 ua1 = 1.033603470734638E-9 lua1 = 1.688934633685681E-16
+ wua1 = 3.424398378187646E-16 pua1 = -2.97233656655428E-22 ub1 = -1.014067449348043E-18
+ lub1 = 1.335471292320971E-25 wub1 = 1.554592007787752E-25 pub1 = -4.950223128976067E-32
+ uc1 = -8.839772191220768E-11 luc1 = 7.867956744515836E-17 wuc1 = 8.252637953539383E-17
+ puc1 = -5.643497257892364E-23 at = 1.278860841856492E5 lat = -0.015875978849476
+ wat = -7.922657276091328E-3 pat = -1.644957070180493E-8 prt = 0
+ njs = 1.2928 xtis = 2 tpb = 1.2287E-3
+ tpbsw = 0 tpbswg = 0 tcj = 7.92E-4
+ tcjsw = 1E-5 tcjswg = 0 tvoff = 0
+ tvfbsdoff = 0 saref = 2.75E-6 sbref = 2.74E-6
+ wlod = 0 ku0 = -2.7E-8 kvsat = 0.2
+ kvth0 = 9.8E-9 tku0 = 0 llodku0 = 0
+ wlodku0 = 1 llodvth = 0 wlodvth = 1
+ lku0 = 0 wku0 = 0 pku0 = 0
+ lkvth0 = 0 wkvth0 = 2E-7 pkvth0 = 0
+ stk2 = 0 lodk2 = 1 steta0 = 0
+ lodeta0 = 1

.model nshort_model.38 nmos
+ level = 54 lmin = 2.5E-7 lmax = 5E-7 wmin = 5.5E-7
+ wmax = 1E-6 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 4.148E-9
+ toxm = 4.148E-9 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 9.999999999999999E22 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {2.1859E-8+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {1.1932E-8-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = 0 dwb = 0 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = 0.629734017174034 lvth0 = -1.803834197187924E-8
+ wvth0 = -8.306347668951688E-9 pvth0 = -1.781089582237517E-15 k1 = 0.177811864220334
+ lk1 = 2.310450597874676E-7 wk1 = 7.161464691227428E-8 pk1 = -7.943621088826815E-14
+ k2 = 0.085399813860113 lk2 = -7.150051800491712E-8 wk2 = -2.550719953689193E-8
+ pk2 = 2.545889332162967E-14 k3 = 2 k3b = 0.54
+ w0 = 0 lpe0 = 1.0325E-7 lpeb = -7.082E-8
+ vbm = -3 dvtp0 = 0 dvtp1 = 0
+ dvt0 = 0 dvt1 = 0.53 dvt2 = -0.032
+ dvt0w = -3.58 dvt1w = 1.6706E6 dvt2w = 0.068
+ vfbsdoff = 0 u0 = 0.018684783930797 lu0 = 1.920004809008676E-9
+ wu0 = 6.541354869874765E-10 pu0 = -6.200987437699484E-16 ua = -2.01231037339091E-9
+ lua = 2.327016480756184E-16 wua = 2.335019899524815E-16 pua = -9.387675945084795E-23
+ ub = 2.511461576438438E-18 lub = -2.265090320778557E-25 wub = -3.763247903905083E-25
+ pub = 1.456027350846167E-31 uc = 9.097622043340024E-11 luc = 6.99631027229822E-18
+ wuc = -2.584110291252102E-17 puc = -5.043499386821734E-25 ud = 0
+ up = 0 lp = 1 eu = 1.67
+ vsat = 4.903866393305725E3 lvsat = 0.031642311110751 wvsat = 0.082307916730562
+ pvsat = -1.494797398457745E-8 a0 = 1.67662360993664 la0 = -2.227859566296791E-8
+ wa0 = -1.689019789574298E-7 pa0 = 2.130462001777428E-14 ags = 2.297500718979647
+ lags = -6.947547928718143E-8 wags = -1.283640403856454E-6 pags = 1.301936499672723E-13
+ b0 = 0 b1 = 0 keta = 0.031694965602808
+ lketa = -4.329897622663901E-8 wketa = -1.60194429333717E-8 pketa = 2.019383755550638E-14
+ a1 = 0 a2 = 0.42385546 rdsw = 65.968
+ rdswmin = 0 rdw = 0 rdwmin = 0
+ rsw = 0 rswmin = 0 prwb = 0
+ prwg = 0.021507 wr = 1 voff = -0.109864841842599
+ lvoff = -1.790461047849649E-8 wvoff = -5.440038436623488E-9 pvoff = 3.514031957455247E-15
+ voffl = 5.8197729E-9 minv = 0 nfactor = 4.714663109597307
+ lnfactor = -6.792621039772253E-7 wnfactor = -8.158414590909653E-7 pnfactor = 3.149792378909037E-13
+ eta0 = 1.232158358211346 leta0 = -3.533683120453174E-7 weta0 = -2.864635283639359E-7
+ peta0 = 1.36395598541091E-13 etab = 0.066426103903855 letab = -3.160924976506588E-8
+ wetab = -2.603300545166505E-8 petab = 1.223516742733478E-14 dsub = 0.097675040093113
+ ldsub = 1.043267293551407E-7 wdsub = 8.058997027729918E-8 pdsub = -3.993363395726089E-14
+ cit = 0 cdsc = 0 cdscb = 0
+ cdscd = 0.010478104286239 lcdscd = -2.417868262432559E-9 wcdscd = -1.960082584226952E-9
+ pcdscd = 9.332658813234838E-16 pclm = 0.939791554400215 lpclm = -1.835858418318944E-7
+ wpclm = -1.94428020640933E-7 ppclm = 6.788799954988178E-14 pdiblc1 = -0.01679926924381
+ lpdiblc1 = 1.341033428627282E-7 wpdiblc1 = -3.387701972515028E-8 ppdiblc1 = -3.975180963093108E-14
+ pdiblc2 = -6.321902690714234E-3 lpdiblc2 = 4.610010848751184E-9 wpdiblc2 = 1.698884552100347E-9
+ ppdiblc2 = -1.607719299658195E-15 pdiblcb = 0.200288832728148 lpdiblcb = -6.998152737554013E-8
+ wpdiblcb = -1.477138813998771E-7 ppdiblcb = 3.467539576626017E-14 drout = 1.753332791971738
+ ldrout = -3.586888086695696E-7 wdrout = -2.907765743253805E-7 pdrout = 1.384491437662194E-13
+ pscbe1 = 1.368678863823744E9 lpscbe1 = -76.28576380166673 wpscbe1 = -536.3955647875989
+ ppscbe1 = 6.94169182969368E-5 pscbe2 = 1E-12 pvag = 0
+ delta = 0.01 fprout = 0 pdits = 0
+ pditsl = 0 pditsd = 0 lambda = 0
+ vtl = 0 lc = 5E-9 xn = 3
+ alpha0 = -5.877019471077723E-6 lalpha0 = 7.394364802538612E-13 walpha0 = 5.656042386662573E-12
+ palpha0 = -7.105693969681459E-19 alpha1 = 0.85 beta0 = 6.607764143963018
+ lbeta0 = 1.225664613657542E-6 wbeta0 = 6.537283001995075E-6 pbeta0 = -9.826266808525891E-13
+ aigbacc = 1 bigbacc = 0 cigbacc = 0
+ nigbacc = 0 aigbinv = 0.35 bigbinv = 0.03
+ cigbinv = 6E-3 eigbinv = 1.1 nigbinv = 0
+ aigc = 0.43 bigc = 0.054 cigc = 0.075
+ aigsd = 0.43 bigsd = 0.054 cigsd = 0.075
+ dlcig = 0 nigc = 0 poxedge = 1
+ pigcd = 1 ntox = 1 toxref = 4.148E-9
+ agidl = 0 bgidl = 2.3E9 cgidl = 0.5
+ egidl = 0.8 noia = 2.5E42 noib = 0
+ noic = 0 em = 4.1E7 af = 1
+ ef = 0.84 kf = 0 lintnoi = -1E-7
+ tnoia = 1.5E7 tnoib = 9.9E6 ntnoi = 1
+ rnoia = 0.94 rnoib = 0.26 xpart = 0
+ cgso = {2.449068E-10/sw_func_tox_lv_ratio} cgdo = {2.449068E-10/sw_func_tox_lv_ratio} cgbo = {1E-13/sw_func_tox_lv_ratio}
+ ckappas = 0.6 cf = 1.4067E-12 clc = 1E-7
+ cle = 0.6 dlc = 9.87908E-9 dwc = 0
+ vfbcv = -1 noff = 3.4037 voffcv = -0.17287
+ acde = 0.4 moin = 6.9 cgsl = {0/sw_func_tox_lv_ratio}
+ cgdl = {0/sw_func_tox_lv_ratio} ijthsrev = 0.1 ijthsfwd = 0.1
+ xjbvs = 1 bvs = 11.7 jss = 2.75E-3
+ jsws = 6E-10 cjs = {sw_nsd_pw_cj} mjs = 0.44
+ mjsws = 9E-4 cjsws = {3.67354204E-11*sw_func_nsd_pw_cj} cjswgs = {2.38232788E-10*sw_func_nsd_pw_cj}
+ mjswgs = 0.8 pbs = 0.729 pbsws = 0.2
+ pbswgs = 0.95578 xrcrg1 = 12 xrcrg2 = 1
+ rbpb = 50 rbpd = 50 rbps = 50
+ rbdb = 50 rbsb = 50 gbmin = 1E-12
+ tnom = 30 ute = -0.929713307571486 lute = -9.587031469188749E-8
+ wute = -2.02751718244245E-7 pute = 5.333601277295477E-14 kt1 = -0.303433900757681
+ lkt1 = 1.994175135536696E-8 wkt1 = 5.464593740513412E-9 pkt1 = -6.795871573135192E-15
+ kt1l = 0 kt2 = -0.047118552144382 lkt2 = 5.324519836093592E-9
+ wkt2 = 3.834897770622467E-9 pkt2 = -2.014638474541086E-15 ua1 = 3.189447151101728E-9
+ lua1 = -8.575813232266965E-16 wua1 = -1.037604234607266E-15 pua1 = 3.598550078132124E-22
+ ub1 = -2.857482412753743E-18 lub1 = 1.011263356248233E-24 wub1 = 8.823560100278814E-25
+ pub1 = -3.956039704583931E-31 uc1 = -7.337056955241399E-11 luc1 = 7.152459922917563E-17
+ wuc1 = 1.42445174437161E-17 puc1 = -2.392351989004058E-23 at = 1.531586071897429E5
+ lat = -0.027909136862554 wat = -0.080004485434936 pat = 1.787118263043468E-8
+ prt = 0 njs = 1.2928 xtis = 2
+ tpb = 1.2287E-3 tpbsw = 0 tpbswg = 0
+ tcj = 7.92E-4 tcjsw = 1E-5 tcjswg = 0
+ tvoff = 0 tvfbsdoff = 0 saref = 1.75E-6
+ sbref = 1.74E-6 wlod = 0 ku0 = -2.7E-8
+ kvsat = 0.2 kvth0 = 9.8E-9 tku0 = 0
+ llodku0 = 0 wlodku0 = 1 llodvth = 0
+ wlodvth = 1 lku0 = 0 wku0 = 0
+ pku0 = 0 lkvth0 = 0 wkvth0 = 2E-7
+ pkvth0 = 0 stk2 = 0 lodk2 = 1
+ steta0 = 0 lodeta0 = 1

.model nshort_model.39 nmos
+ level = 54 lmin = 1.8E-7 lmax = 2.5E-7 wmin = 5.5E-7
+ wmax = 1E-6 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 4.148E-9
+ toxm = 4.148E-9 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 9.999999999999999E22 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {2.1859E-8+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {1.1932E-8-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = 0 dwb = 0 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = 0.621261040746794 lvth0 = -1.612229697452869E-8
+ wvth0 = -4.016632217414285E-9 pvth0 = -2.75114867558638E-15 k1 = 1.568401017801571
+ lk1 = -8.341720904677905E-8 wk1 = -6.324156109411419E-7 pk1 = 7.977037550167196E-14
+ k2 = -0.372944893267147 lk2 = 3.214772068601298E-8 wk2 = 2.065444754769111E-7
+ pk2 = -2.701634425929168E-14 k3 = 2 k3b = 0.54
+ w0 = 0 lpe0 = 1.0325E-7 lpeb = -7.082E-8
+ vbm = -3 dvtp0 = 0 dvtp1 = 0
+ dvt0 = 0 dvt1 = 0.53 dvt2 = -0.032
+ dvt0w = -3.58 dvt1w = 1.6706E6 dvt2w = 0.068
+ vfbsdoff = 0 u0 = 0.024624633295691 lu0 = 5.767910330288167E-10
+ wu0 = -2.353103329171248E-9 pu0 = 5.994621316092093E-17 ua = -7.260331848850542E-10
+ lua = -5.817193022434168E-17 wua = -4.177169975986398E-16 pua = 5.338729751801239E-23
+ ub = 1.131725908750084E-18 lub = 8.549887287051786E-26 wub = 3.222105429180885E-25
+ pub = -1.236125104845611E-32 uc = 6.820031183327979E-11 luc = 1.214676313949506E-17
+ wuc = -1.431007035463473E-17 puc = -3.111931517192347E-24 ud = 0
+ up = 0 lp = 1 eu = 1.67
+ vsat = 7.753122894440708E4 lvsat = 0.015218649852896 wvsat = 0.045537990363465
+ pvsat = -6.63296991562763E-9 a0 = 1.67662360993664 la0 = -2.22785956629681E-8
+ wa0 = -1.689019789574305E-7 pa0 = 2.130462001777446E-14 ags = 2.924021433000002
+ lags = -2.111543674728882E-7 wags = -1.600836563992108E-6 pags = 2.019231208357085E-13
+ b0 = 0 b1 = 0 keta = -0.38601732580332
+ lketa = 5.11608105027772E-8 wketa = 1.954607713843063E-7 pketa = -2.762945218943604E-14
+ a1 = 0 a2 = 0.42385546 rdsw = 65.968
+ rdswmin = 0 rdw = 0 rdwmin = 0
+ rsw = 0 rswmin = 0 prwb = 0
+ prwg = 0.021507 wr = 1 voff = -0.105890915176759
+ lvoff = -1.880325835900282E-8 wvoff = -7.451965976858132E-9 pvoff = 3.969001203693748E-15
+ voffl = 5.8197729E-9 minv = 0 nfactor = 6.362854041802729
+ lnfactor = -1.051977408622431E-6 wnfactor = -1.65029086062979E-6 pnfactor = 5.036782877572874E-13
+ eta0 = -0.748205051907289 leta0 = 9.44631480652703E-8 weta0 = 7.161588196377473E-7
+ peta0 = -9.033340874661768E-14 etab = -0.110381846046637 letab = 8.3733928049386E-9
+ wetab = 6.348167706517028E-8 petab = -8.007324818292297E-15 dsub = 0.685664590572337
+ ldsub = -2.863887563202906E-8 wdsub = -2.170985553184241E-7 pdsub = 2.738445846685357E-14
+ cit = 0 cdsc = 0 cdscb = 0
+ cdscd = -3.072227435596798E-3 lcdscd = 6.463495518164379E-10 wcdscd = 4.900206460567379E-9
+ pcdscd = -6.180924421101269E-16 pclm = 0.397941715007052 lpclm = -6.105408655088194E-8
+ wpclm = 7.990079974671711E-8 ppclm = 5.852377422700131E-15 pdiblc1 = 0.852773842006099
+ lpdiblc1 = -6.25384422228814E-8 wpdiblc1 = -4.741262336349769E-7 ppdiblc1 = 5.980438660578147E-14
+ pdiblc2 = 0.021200877060382 lpdiblc2 = -1.613880473042784E-9 wpdiblc2 = -1.223540342584432E-8
+ ppdiblc2 = 1.5433248465223E-15 pdiblcb = -0.116596966530078 lpdiblcb = 1.677759725518053E-9
+ wpdiblcb = 1.271969482017651E-8 ppdiblcb = -1.604411425837855E-15 drout = -0.256848118894546
+ ldrout = 9.588546179008854E-8 wdrout = 7.269414579108348E-7 pdrout = -9.169354117154945E-14
+ pscbe1 = 1.333952617642992E9 lpscbe1 = -68.43290939533645 wpscbe1 = -518.8142914187162
+ ppscbe1 = 6.544115946239114E-5 pscbe2 = 1E-12 pvag = 0
+ delta = 0.01 fprout = 0 pdits = 0
+ pditsl = 0 pditsd = 0 lambda = 0
+ vtl = 0 lc = 5E-9 xn = 3
+ alpha0 = -5.911016719125336E-6 lalpha0 = 7.471244819383567E-13 walpha0 = 5.673254581398614E-12
+ palpha0 = -7.144616938369757E-19 alpha1 = 0.85 beta0 = 9.607118556871509
+ lbeta0 = 5.474026041400681E-7 wbeta0 = 5.018763851118943E-6 pbeta0 = -6.392348341500643E-13
+ aigbacc = 1 bigbacc = 0 cigbacc = 0
+ nigbacc = 0 aigbinv = 0.35 bigbinv = 0.03
+ cigbinv = 6E-3 eigbinv = 1.1 nigbinv = 0
+ aigc = 0.43 bigc = 0.054 cigc = 0.075
+ aigsd = 0.43 bigsd = 0.054 cigsd = 0.075
+ dlcig = 0 nigc = 0 poxedge = 1
+ pigcd = 1 ntox = 1 toxref = 4.148E-9
+ agidl = 0 bgidl = 2.3E9 cgidl = 0.5
+ egidl = 0.8 noia = 2.5E42 noib = 0
+ noic = 0 em = 4.1E7 af = 1
+ ef = 0.84 kf = 0 lintnoi = -1E-7
+ tnoia = 1.5E7 tnoib = 9.9E6 ntnoi = 1
+ rnoia = 0.94 rnoib = 0.26 xpart = 0
+ cgso = {2.449068E-10/sw_func_tox_lv_ratio} cgdo = {2.449068E-10/sw_func_tox_lv_ratio} cgbo = {1E-13/sw_func_tox_lv_ratio}
+ ckappas = 0.6 cf = 1.4067E-12 clc = 1E-7
+ cle = 0.6 dlc = 9.87908E-9 dwc = 0
+ vfbcv = -1 noff = 3.4037 voffcv = -0.17287
+ acde = 0.4 moin = 6.9 cgsl = {0/sw_func_tox_lv_ratio}
+ cgdl = {0/sw_func_tox_lv_ratio} ijthsrev = 0.1 ijthsfwd = 0.1
+ xjbvs = 1 bvs = 11.7 jss = 2.75E-3
+ jsws = 6E-10 cjs = {sw_nsd_pw_cj} mjs = 0.44
+ mjsws = 9E-4 cjsws = {3.67354204E-11*sw_func_nsd_pw_cj} cjswgs = {2.38232788E-10*sw_func_nsd_pw_cj}
+ mjswgs = 0.8 pbs = 0.729 pbsws = 0.2
+ pbswgs = 0.95578 xrcrg1 = 12 xrcrg2 = 1
+ rbpb = 50 rbpd = 50 rbps = 50
+ rbdb = 50 rbsb = 50 gbmin = 1E-12
+ tnom = 30 ute = -1.306507640787219 lute = -1.066355135581445E-8
+ wute = -1.198752963511675E-8 pute = 1.019736221764095E-14 kt1 = -0.182817533257321
+ lkt1 = -7.333951525694416E-9 wkt1 = -5.560130203030283E-8 pkt1 = 7.013325832894108E-15
+ kt1l = 0 kt2 = -0.016880072219243 lkt2 = -1.513489060257432E-9
+ wkt2 = -1.147430032283539E-8 pkt2 = 1.447322345521098E-15 ua1 = -1.333244946914602E-9
+ lua1 = 1.651621770503242E-16 wua1 = 1.252153366160638E-15 pua1 = -1.579416169940382E-22
+ ub1 = 2.758105595066333E-18 lub1 = -2.58623253488167E-25 wub1 = -1.960715117747282E-24
+ pub1 = 2.473167620921713E-31 uc1 = 3.636738728287094E-10 luc1 = -2.730688279312209E-17
+ wuc1 = -2.070232169338839E-16 puc1 = 2.611308049117238E-23 at = -8.517354882322786E4
+ lat = 0.025986343569596 wat = 0.040658795175622 pat = -9.415128993714486E-9
+ prt = 0 njs = 1.2928 xtis = 2
+ tpb = 1.2287E-3 tpbsw = 0 tpbswg = 0
+ tcj = 7.92E-4 tcjsw = 1E-5 tcjswg = 0
+ tvoff = 0 tvfbsdoff = 0 saref = 1.75E-6
+ sbref = 1.74E-6 wlod = 0 ku0 = -2.7E-8
+ kvsat = 0.2 kvth0 = 9.8E-9 tku0 = 0
+ llodku0 = 0 wlodku0 = 1 llodvth = 0
+ wlodvth = 1 lku0 = 0 wku0 = 0
+ pku0 = 0 lkvth0 = 0 wkvth0 = 2E-7
+ pkvth0 = 0 stk2 = 0 lodk2 = 1
+ steta0 = 0 lodeta0 = 1

.model nshort_model.40 nmos
+ level = 54 lmin = 1.5E-7 lmax = 1.8E-7 wmin = 5.5E-7
+ wmax = 1E-6 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 4.148E-9
+ toxm = 4.148E-9 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 9.999999999999999E22 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {2.1859E-8+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {1.1932E-8-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = 0 dwb = 0 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = 0.561743750427059 lvth0 = -6.829505333166525E-9
+ wvth0 = 2.611590056024244E-8 pvth0 = -7.455921813358589E-15 k1 = 1.568401017801568
+ lk1 = -8.34172090467785E-8 wk1 = -6.324156109411386E-7 pk1 = 7.977037550167143E-14
+ k2 = -0.35166619774707 lk2 = 2.88253502822903E-8 wk2 = 1.957714549516151E-7
+ pk2 = -2.533428792655407E-14 k3 = 2 k3b = 0.54
+ w0 = 0 lpe0 = 1.0325E-7 lpeb = -7.082E-8
+ vbm = -3 dvtp0 = 0 dvtp1 = 0
+ dvt0 = 0 dvt1 = 0.53 dvt2 = -0.032
+ dvt0w = -3.58 dvt1w = 1.6706E6 dvt2w = 0.068
+ vfbsdoff = 0 u0 = 0.033073526744731 lu0 = -7.423853945304192E-10
+ wu0 = -6.630626002339119E-9 pu0 = 7.278214932586596E-16 ua = -7.595255951297886E-10
+ lua = -5.294255925836984E-17 wua = -4.007603931551177E-16 pua = 5.073976112661863E-23
+ ub = 2.951933331337695E-18 lub = -1.987010332626215E-25 wub = -5.993277114044132E-25
+ pub = 1.31524045828442E-31 uc = 4.498456474434723E-10 luc = -4.744181298133794E-17
+ wuc = -2.075302341580341E-16 puc = 2.705669197841522E-23 ud = 0
+ up = 0 lp = 1 eu = 1.67
+ vsat = 1.654122069777363E5 lvsat = 1.49726546668362E-3 wvsat = 1.045433042794898E-3
+ pvsat = 3.139200141924857E-10 a0 = 1.67662360993664 la0 = -2.227859566296807E-8
+ wa0 = -1.689019789574304E-7 pa0 = 2.130462001777443E-14 ags = 2.924021433000002
+ lags = -2.111543674728881E-7 wags = -1.600836563992107E-6 pags = 2.019231208357084E-13
+ b0 = 0 b1 = 0 keta = -0.431400461998999
+ lketa = 5.824675185582569E-8 wketa = 2.184374363437266E-7 pketa = -3.121693674954008E-14
+ a1 = 0 a2 = 0.42385546 rdsw = 65.968
+ rdswmin = 0 rdw = 0 rdwmin = 0
+ rsw = 0 rswmin = 0 prwb = 0
+ prwg = 0.021507 wr = 1 voff = -0.305321273701378
+ lvoff = 1.233500009959698E-8 wvoff = 9.351603479770085E-8 pvoff = -1.179573856524279E-14
+ voffl = 5.8197729E-9 minv = 0 nfactor = -15.04415574837766
+ lnfactor = 2.290427471977174E-6 wnfactor = 9.187692869962315E-6 pnfactor = -1.188521140002441E-12
+ eta0 = -0.748205060282676 leta0 = 9.446314937296974E-8 weta0 = 7.161588238780545E-7
+ peta0 = -9.033340940868227E-14 etab = -0.110381846046638 letab = 8.373392804938716E-9
+ wetab = 6.348167706517098E-8 petab = -8.007324818292406E-15 dsub = 0.685630677113776
+ ldsub = -2.863358052026326E-8 wdsub = -2.170813855447961E-7 pdsub = 2.738177764707839E-14
+ cit = 0 cdsc = 0 cdscb = 0
+ cdscd = -3.072227435596797E-3 lcdscd = 6.463495518164378E-10 wcdscd = 4.900206460567378E-9
+ pcdscd = -6.180924421101268E-16 pclm = -0.349733339964259 lpclm = 5.568490583211858E-8
+ wpclm = 4.584352219277013E-7 ppclm = -5.325047311895002E-14 pdiblc1 = 0.852773842006098
+ lpdiblc1 = -6.253844222288121E-8 wpdiblc1 = -4.741262336349758E-7 ppdiblc1 = 5.98043866057813E-14
+ pdiblc2 = 0.021200877060382 lpdiblc2 = -1.61388047304278E-9 wpdiblc2 = -1.22354034258443E-8
+ ppdiblc2 = 1.543324846522296E-15 pdiblcb = -0.116596966530076 lpdiblcb = 1.677759725517667E-9
+ wpdiblcb = 1.271969482017414E-8 ppdiblcb = -1.604411425837486E-15 drout = -0.256846256246345
+ ldrout = 9.588517096364904E-8 wdrout = 7.269396766938879E-7 pdrout = -9.169326305946023E-14
+ pscbe1 = 1.333952617642994E9 lpscbe1 = -68.43290939533665 wpscbe1 = -518.8142914187174
+ ppscbe1 = 6.544115946239133E-5 pscbe2 = 1E-12 pvag = 0
+ delta = 0.01 fprout = 0 pdits = 0
+ pditsl = 0 pditsd = 0 lambda = 0
+ vtl = 0 lc = 5E-9 xn = 3
+ alpha0 = -5.986070150633222E-6 lalpha0 = 7.588430245202721E-13 walpha0 = 5.71125278280928E-12
+ palpha0 = -7.203945810124312E-19 alpha1 = 0.85 beta0 = 10.014535571191939
+ lbeta0 = 4.837901411921336E-7 wbeta0 = 4.812495950274766E-6 pbeta0 = -6.070289891838577E-13
+ aigbacc = 1 bigbacc = 0 cigbacc = 0
+ nigbacc = 0 aigbinv = 0.35 bigbinv = 0.03
+ cigbinv = 6E-3 eigbinv = 1.1 nigbinv = 0
+ aigc = 0.43 bigc = 0.054 cigc = 0.075
+ aigsd = 0.43 bigsd = 0.054 cigsd = 0.075
+ dlcig = 0 nigc = 0 poxedge = 1
+ pigcd = 1 ntox = 1 toxref = 4.148E-9
+ agidl = 0 bgidl = 2.3E9 cgidl = 0.5
+ egidl = 0.8 noia = 2.5E42 noib = 0
+ noic = 0 em = 4.1E7 af = 1
+ ef = 0.84 kf = 0 lintnoi = -1E-7
+ tnoia = 1.5E7 tnoib = 9.9E6 ntnoi = 1
+ rnoia = 0.94 rnoib = 0.26 xpart = 0
+ cgso = {2.449068E-10/sw_func_tox_lv_ratio} cgdo = {2.449068E-10/sw_func_tox_lv_ratio} cgbo = {1E-13/sw_func_tox_lv_ratio}
+ ckappas = 0.6 cf = 1.4067E-12 clc = 1E-7
+ cle = 0.6 dlc = 9.87908E-9 dwc = 0
+ vfbcv = -1 noff = 3.4037 voffcv = -0.17287
+ acde = 0.4 moin = 6.9 cgsl = {0/sw_func_tox_lv_ratio}
+ cgdl = {0/sw_func_tox_lv_ratio} ijthsrev = 0.1 ijthsfwd = 0.1
+ xjbvs = 1 bvs = 11.7 jss = 2.75E-3
+ jsws = 6E-10 cjs = {sw_nsd_pw_cj} mjs = 0.44
+ mjsws = 9E-4 cjsws = {3.67354204E-11*sw_func_nsd_pw_cj} cjswgs = {2.38232788E-10*sw_func_nsd_pw_cj}
+ mjswgs = 0.8 pbs = 0.729 pbsws = 0.2
+ pbswgs = 0.95578 xrcrg1 = 12 xrcrg2 = 1
+ rbpb = 50 rbpd = 50 rbps = 50
+ rbdb = 50 rbsb = 50 gbmin = 1E-12
+ tnom = 30 ute = -1.306507640787218 lute = -1.066355135581462E-8
+ wute = -1.198752963511782E-8 pute = 1.019736221764112E-14 kt1 = -0.361516179704722
+ lkt1 = 2.056734033601708E-8 wkt1 = 3.487060609037792E-8 pkt1 = -7.112596013436501E-15
+ kt1l = 0 kt2 = -0.016880072219241 lkt2 = -1.51348906025779E-9
+ wkt2 = -1.147430032283757E-8 pkt2 = 1.44732234552144E-15 ua1 = -1.333244946914601E-9
+ lua1 = 1.651621770503241E-16 wua1 = 1.252153366160637E-15 pua1 = -1.579416169940381E-22
+ ub1 = 2.758105595066328E-18 lub1 = -2.586232534881663E-25 wub1 = -1.960715117747278E-24
+ pub1 = 2.473167620921706E-31 uc1 = 3.636738728287096E-10 luc1 = -2.730688279312211E-17
+ wuc1 = -2.070232169338841E-16 puc1 = 2.61130804911724E-23 at = 3.132074202674847E5
+ lat = -0.036215267420352 wat = -0.161034318617564 pat = 2.20764270214984E-8
+ prt = 0 njs = 1.2928 xtis = 2
+ tpb = 1.2287E-3 tpbsw = 0 tpbswg = 0
+ tcj = 7.92E-4 tcjsw = 1E-5 tcjswg = 0
+ tvoff = 0 tvfbsdoff = 0 saref = 1.75E-6
+ sbref = 1.74E-6 wlod = 0 ku0 = -2.7E-8
+ kvsat = 0.2 kvth0 = 9.8E-9 tku0 = 0
+ llodku0 = 0 wlodku0 = 1 llodvth = 0
+ wlodvth = 1 lku0 = 0 wku0 = 0
+ pku0 = 0 lkvth0 = 0 wkvth0 = 2E-7
+ pkvth0 = 0 stk2 = 0 lodk2 = 1
+ steta0 = 0 lodeta0 = 1

.model nshort_model.41 nmos
+ level = 54 lmin = 8E-6 lmax = 2.02E-5 wmin = 4.2E-7
+ wmax = 5.5E-7 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 4.148E-9
+ toxm = 4.148E-9 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 9.999999999999999E22 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {2.1859E-8+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {1.1932E-8-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = 0 dwb = 0 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = 0.647883369553665 lvth0 = -7.97909620444532E-7
+ wvth0 = -6.501808598696865E-8 pvth0 = 4.039672784578986E-13 k1 = 0.341104073284211
+ lk1 = -6.552377723129526E-7 wk1 = 8.111562450940306E-8 pk1 = 3.317350898421464E-13
+ k2 = 0.027661713114934 lk2 = 4.935418965694249E-7 wk2 = -2.092161565234127E-8
+ pk2 = -2.498713784789616E-13 k3 = 2 k3b = 0.54
+ w0 = 0 lpe0 = 1.0325E-7 lpeb = -7.082E-8
+ vbm = -3 dvtp0 = 0 dvtp1 = 0
+ dvt0 = 0 dvt1 = 0.53 dvt2 = -0.032
+ dvt0w = -3.58 dvt1w = 1.6706E6 dvt2w = 0.068
+ vfbsdoff = 0 u0 = 0.039805665304804 lu0 = -6.857804440511436E-8
+ wu0 = -6.25742544164686E-9 pu0 = 3.471982947751011E-14 ua = 3.031964223296942E-10
+ lua = -5.104678065069638E-15 wua = -5.438404098418022E-16 pua = 2.584406620139586E-21
+ ub = 9.599749736472269E-19 lub = 2.376634311820368E-24 wub = 2.550547441134748E-25
+ pub = -1.20324717265704E-30 uc = -8.077411491515575E-11 luc = 8.545737476978952E-16
+ wuc = 5.421881012347488E-17 puc = -4.326553061319858E-22 ud = 0
+ up = 0 lp = 1 eu = 1.67
+ vsat = 8E4 a0 = 0.860783192981373 la0 = 6.710225595792974E-6
+ wa0 = 2.324932034910048E-7 pa0 = -3.397266435089259E-12 ags = 0.553423993594853
+ lags = -1.355111996034707E-6 wags = -8.729010150518953E-8 pags = 6.860688115764437E-13
+ b0 = 4.899303586829902E-8 lb0 = -6.180248442494087E-13 wb0 = -1.367925151747417E-14
+ pb0 = 3.128948541962792E-19 b1 = -4.578338796966269E-9 lb1 = 1.831668682104781E-14
+ wb1 = 3.313736588605676E-15 pb1 = -9.273408837133729E-21 keta = -0.023060366272357
+ lketa = 1.49062319563818E-7 wketa = 7.936459556301426E-9 pketa = -7.546756927340891E-14
+ a1 = 0 a2 = 0.42385546 rdsw = 65.968
+ rdswmin = 0 rdw = 0 rdwmin = 0
+ rsw = 0 rswmin = 0 prwb = 0
+ prwg = 0.021507 wr = 1 voff = -0.165762140220576
+ lvoff = 3.768045323177115E-7 wvoff = 2.408246282745343E-8 pvoff = -1.907693522308756E-13
+ voffl = 5.8197729E-9 minv = 0 nfactor = 0.986789554983682
+ lnfactor = 9.592624906700605E-6 wnfactor = 9.498915765237517E-7 pnfactor = -4.856573323014196E-12
+ eta0 = 0.08 etab = -0.07 dsub = 0.56
+ cit = 0 cdsc = 0 cdscb = 0
+ cdscd = 5.4E-3 pclm = 0.300893230860127 lpclm = -2.561722779571456E-6
+ wpclm = -1.23542037956327E-7 ppclm = 1.296954132286996E-12 pdiblc1 = 0.39
+ pdiblc2 = 6.5828309153609E-3 lpdiblc2 = -6.448342862049019E-8 wpdiblc2 = -2.535289849255748E-9
+ ppdiblc2 = 3.264679920883902E-14 pdiblcb = -0.025 drout = 0.56
+ pscbe1 = 2.820123968488849E9 lpscbe1 = -1.683214049179674E4 wpscbe1 = -1.086038052977252E3
+ ppscbe1 = 8.521809752467836E-3 pscbe2 = 1E-12 pvag = 0
+ delta = 0.01 fprout = 0 pdits = 0
+ pditsl = 0 pditsd = 0 lambda = 0
+ vtl = 0 lc = 5E-9 xn = 3
+ alpha0 = 3E-8 alpha1 = 0.85 beta0 = 13.86
+ aigbacc = 1 bigbacc = 0 cigbacc = 0
+ nigbacc = 0 aigbinv = 0.35 bigbinv = 0.03
+ cigbinv = 6E-3 eigbinv = 1.1 nigbinv = 0
+ aigc = 0.43 bigc = 0.054 cigc = 0.075
+ aigsd = 0.43 bigsd = 0.054 cigsd = 0.075
+ dlcig = 0 nigc = 0 poxedge = 1
+ pigcd = 1 ntox = 1 toxref = 4.148E-9
+ agidl = 0 bgidl = 2.3E9 cgidl = 0.5
+ egidl = 0.8 noia = 2.5E42 noib = 0
+ noic = 0 em = 4.1E7 af = 1
+ ef = 0.84 kf = 0 lintnoi = -1E-7
+ tnoia = 1.5E7 tnoib = 9.9E6 ntnoi = 1
+ rnoia = 0.94 rnoib = 0.26 xpart = 0
+ cgso = {2.449068E-10/sw_func_tox_lv_ratio} cgdo = {2.449068E-10/sw_func_tox_lv_ratio} cgbo = {1E-13/sw_func_tox_lv_ratio}
+ ckappas = 0.6 cf = 1.4067E-12 clc = 1E-7
+ cle = 0.6 dlc = 9.87908E-9 dwc = 0
+ vfbcv = -1 noff = 3.4037 voffcv = -0.17287
+ acde = 0.4 moin = 6.9 cgsl = {0/sw_func_tox_lv_ratio}
+ cgdl = {0/sw_func_tox_lv_ratio} ijthsrev = 0.1 ijthsfwd = 0.1
+ xjbvs = 1 bvs = 11.7 jss = 2.75E-3
+ jsws = 6E-10 cjs = {sw_nsd_pw_cj} mjs = 0.44
+ mjsws = 9E-4 cjsws = {3.67354204E-11*sw_func_nsd_pw_cj} cjswgs = {2.38232788E-10*sw_func_nsd_pw_cj}
+ mjswgs = 0.8 pbs = 0.729 pbsws = 0.2
+ pbswgs = 0.95578 xrcrg1 = 12 xrcrg2 = 1
+ rbpb = 50 rbpd = 50 rbps = 50
+ rbdb = 50 rbsb = 50 gbmin = 1E-12
+ tnom = 30 ute = -1.67377733769147 lute = -4.919294823948998E-7
+ wute = 2.069059798811131E-7 pute = 2.490550422058547E-13 kt1 = -0.327696628520005
+ lkt1 = 4.550347712152836E-7 wkt1 = 1.850796300036506E-8 pkt1 = -2.303759140404162E-13
+ kt1l = 0 kt2 = 2.286629874913983E-3 lkt2 = 6.068376760439134E-8
+ wkt2 = -1.15725680722892E-8 pkt2 = -3.072309923028646E-14 ua1 = 2.361964247265615E-9
+ lua1 = -1.41237566234474E-14 wua1 = -5.588665988341301E-16 pua1 = 7.150603750832199E-21
+ ub1 = -2.593080470692032E-18 lub1 = 1.855996132288832E-23 wub1 = 8.822320630429032E-25
+ pub1 = -9.396574338474542E-30 uc1 = -2.011743423026584E-10 luc1 = 5.401421458447489E-16
+ wuc1 = 9.193864294742451E-17 puc1 = -2.734642458825712E-22 at = 215.40504676935234
+ lat = 0.768639816242036 wat = 0.070770424302112 pat = -3.891485034466503E-7
+ prt = 0 njs = 1.2928 xtis = 2
+ tpb = 1.2287E-3 tpbsw = 0 tpbswg = 0
+ tcj = 7.92E-4 tcjsw = 1E-5 tcjswg = 0
+ tvoff = 0 tvfbsdoff = 0 saref = 3E-6
+ sbref = 3E-6 wlod = 0 ku0 = -2.7E-8
+ kvsat = 0.2 kvth0 = 9.8E-9 tku0 = 0
+ llodku0 = 0 wlodku0 = 1 llodvth = 0
+ wlodvth = 1 lku0 = 0 wku0 = 0
+ pku0 = 0 lkvth0 = 0 wkvth0 = 2E-7
+ pkvth0 = 0 stk2 = 0 lodk2 = 1
+ steta0 = 0 lodeta0 = 1

.model nshort_model.42 nmos
+ level = 54 lmin = 4E-6 lmax = 8E-6 wmin = 4.2E-7
+ wmax = 5.5E-7 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 4.148E-9
+ toxm = 4.148E-9 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 9.999999999999999E22 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {2.1859E-8+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {1.1932E-8-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = 0 dwb = 0 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = 0.518512321511687 lvth0 = 2.33971453200822E-7
+ wvth0 = -3.320584705516613E-9 pvth0 = -8.814038262313726E-14 k1 = -0.05609894092055
+ lk1 = 2.512907488594155E-6 wk1 = 2.496208730477575E-7 pk1 = -1.01228568921357E-12
+ k2 = 0.224995014655131 lk2 = -1.08041535384419E-6 wk2 = -1.064235050767482E-7
+ pk2 = 4.321033198270697E-13 k3 = 2 k3b = 0.54
+ w0 = 0 lpe0 = 1.0325E-7 lpeb = -7.082E-8
+ vbm = -3 dvtp0 = 0 dvtp1 = 0
+ dvt0 = 0 dvt1 = 0.53 dvt2 = -0.032
+ dvt0w = -3.58 dvt1w = 1.6706E6 dvt2w = 0.068
+ vfbsdoff = 0 u0 = 0.030218433300949 lu0 = 7.891021921189781E-9
+ wu0 = -2.278099994334348E-9 pu0 = 2.980188521484672E-15 ua = -2.397756544095677E-10
+ lua = -7.73858936794851E-16 wua = -3.731722689570105E-16 pua = 1.223134317575327E-21
+ ub = 1.079815624262907E-18 lub = 1.420768984181218E-24 wub = 2.774926887232715E-25
+ pub = -1.382215270425246E-30 uc = -5.687251165149655E-11 luc = 6.639313094489057E-16
+ wuc = 3.365350308835442E-17 puc = -2.686236203381082E-22 ud = 0
+ up = 0 lp = 1 eu = 1.67
+ vsat = 8E4 a0 = 1.998693023956431 la0 = -2.365897971801105E-6
+ wa0 = -2.983165246117898E-7 pa0 = 8.365441463816526E-13 ags = 0.228950201250347
+ lags = 1.232935100140831E-6 wags = 6.683938675535756E-8 pags = -5.432889484000835E-13
+ b0 = -1.73643685675305E-7 lb0 = 1.157755925376507E-12 wb0 = 9.339313191293379E-14
+ pb0 = -5.411290378888013E-19 b1 = -8.558560960275048E-10 lb1 = -1.13743414592871E-14
+ wb1 = 7.362201388866383E-16 pb1 = 1.128521290806248E-20 keta = -0.012318458536868
+ lketa = 6.338340256610455E-8 wketa = -2.60504680473981E-9 pketa = 8.612919107121094E-15
+ a1 = 0 a2 = 0.42385546 rdsw = 65.968
+ rdswmin = 0 rdw = 0 rdwmin = 0
+ rsw = 0 rswmin = 0 prwb = 0
+ prwg = 0.021507 wr = 1 voff = -0.094852486019431
+ lvoff = -1.887805133035858E-7 wvoff = -1.171828868968579E-8 pvoff = 9.47823107720331E-14
+ voffl = 5.8197729E-9 minv = 0 nfactor = 1.841810105518711
+ lnfactor = 2.772864712838334E-6 wnfactor = 5.031605063882827E-7 pnfactor = -1.293385552188155E-12
+ eta0 = 0.08 etab = -0.07 dsub = 0.56
+ cit = 0 cdsc = 0 cdscb = 0
+ cdscd = 5.4E-3 pclm = -1.705472938229716 lpclm = 1.344132665088813E-5
+ wpclm = 5.118070079259765E-7 ppclm = -3.770676265140497E-12 pdiblc1 = 0.39
+ pdiblc2 = -3.367602183070396E-3 lpdiblc2 = 1.488257903149923E-8 wpdiblc2 = 8.729541800811693E-10
+ ppdiblc2 = 5.462181309659771E-15 pdiblcb = -0.025 drout = 0.56
+ pscbe1 = 9.639156659365531E8 lpscbe1 = -2.026770626310478E3 wpscbe1 = -164.49315042404635
+ ppscbe1 = 1.171442279596724E-3 pscbe2 = 1E-12 pvag = 0
+ delta = 0.01 fprout = 0 pdits = 0
+ pditsl = 0 pditsd = 0 lambda = 0
+ vtl = 0 lc = 5E-9 xn = 3
+ alpha0 = 3E-8 alpha1 = 0.85 beta0 = 13.86
+ aigbacc = 1 bigbacc = 0 cigbacc = 0
+ nigbacc = 0 aigbinv = 0.35 bigbinv = 0.03
+ cigbinv = 6E-3 eigbinv = 1.1 nigbinv = 0
+ aigc = 0.43 bigc = 0.054 cigc = 0.075
+ aigsd = 0.43 bigsd = 0.054 cigsd = 0.075
+ dlcig = 0 nigc = 0 poxedge = 1
+ pigcd = 1 ntox = 1 toxref = 4.148E-9
+ agidl = 0 bgidl = 2.3E9 cgidl = 0.5
+ egidl = 0.8 noia = 2.5E42 noib = 0
+ noic = 0 em = 4.1E7 af = 1
+ ef = 0.84 kf = 0 lintnoi = -1E-7
+ tnoia = 1.5E7 tnoib = 9.9E6 ntnoi = 1
+ rnoia = 0.94 rnoib = 0.26 xpart = 0
+ cgso = {2.449068E-10/sw_func_tox_lv_ratio} cgdo = {2.449068E-10/sw_func_tox_lv_ratio} cgbo = {1E-13/sw_func_tox_lv_ratio}
+ ckappas = 0.6 cf = 1.4067E-12 clc = 1E-7
+ cle = 0.6 dlc = 9.87908E-9 dwc = 0
+ vfbcv = -1 noff = 3.4037 voffcv = -0.17287
+ acde = 0.4 moin = 6.9 cgsl = {0/sw_func_tox_lv_ratio}
+ cgdl = {0/sw_func_tox_lv_ratio} ijthsrev = 0.1 ijthsfwd = 0.1
+ xjbvs = 1 bvs = 11.7 jss = 2.75E-3
+ jsws = 6E-10 cjs = {sw_nsd_pw_cj} mjs = 0.44
+ mjsws = 9E-4 cjsws = {3.67354204E-11*sw_func_nsd_pw_cj} cjswgs = {2.38232788E-10*sw_func_nsd_pw_cj}
+ mjswgs = 0.8 pbs = 0.729 pbsws = 0.2
+ pbswgs = 0.95578 xrcrg1 = 12 xrcrg2 = 1
+ rbpb = 50 rbpd = 50 rbps = 50
+ rbdb = 50 rbsb = 50 gbmin = 1E-12
+ tnom = 30 ute = -2.458926124939385 lute = 5.770524024929533E-6
+ wute = 6.216745483770304E-7 pute = -3.059195468642898E-12 kt1 = -0.296504923284307
+ lkt1 = 2.062454881834426E-7 wkt1 = 5.18214554600651E-9 pkt1 = -1.240873817132786E-13
+ kt1l = 0 kt2 = 0.01560490806981 lkt2 = -4.554463056393125E-8
+ wkt2 = -1.285959395314229E-8 pkt2 = -2.045760576908244E-14 ua1 = -1.022982914455386E-9
+ lua1 = 1.28750422912533E-14 wua1 = 1.28539209572015E-15 pua1 = -7.559454416115196E-21
+ ub1 = 8.857179151784749E-19 lub1 = -9.187407719395327E-24 wub1 = -9.686065248102689E-25
+ pub1 = 5.365965952290307E-30 uc1 = -2.425707490704136E-10 luc1 = 8.703255161356848E-16
+ wuc1 = 8.67604688996675E-17 puc1 = -2.321624254459907E-22 at = 5.342471904753853E4
+ lat = 0.344235091305196 wat = 0.043831506391174 pat = -1.742800304961774E-7
+ prt = 0 njs = 1.2928 xtis = 2
+ tpb = 1.2287E-3 tpbsw = 0 tpbswg = 0
+ tcj = 7.92E-4 tcjsw = 1E-5 tcjswg = 0
+ tvoff = 0 tvfbsdoff = 0 saref = 3E-6
+ sbref = 3E-6 wlod = 0 ku0 = -2.7E-8
+ kvsat = 0.2 kvth0 = 9.8E-9 tku0 = 0
+ llodku0 = 0 wlodku0 = 1 llodvth = 0
+ wlodvth = 1 lku0 = 0 wku0 = 0
+ pku0 = 0 lkvth0 = 0 wkvth0 = 2E-7
+ pkvth0 = 0 stk2 = 0 lodk2 = 1
+ steta0 = 0 lodeta0 = 1

.model nshort_model.43 nmos
+ level = 54 lmin = 2E-6 lmax = 4E-6 wmin = 4.2E-7
+ wmax = 5.5E-7 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 4.148E-9
+ toxm = 4.148E-9 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 9.999999999999999E22 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {2.1859E-8+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {1.1932E-8-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = 0 dwb = 0 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = 0.614532311736839 lvth0 = -1.478170866530562E-7
+ wvth0 = -3.994044756595567E-8 pvth0 = 5.746517241131747E-14 k1 = 0.666711467554453
+ lk1 = -3.610849977180101E-7 wk1 = -5.445611371352468E-8 pk1 = 1.967657646194876E-13
+ k2 = -0.090849395294886 lk2 = 1.754249749568312E-7 wk2 = 2.589283866120042E-8
+ pk2 = -9.400445789776231E-14 k3 = 2 k3b = 0.54
+ w0 = 0 lpe0 = 1.0325E-7 lpeb = -7.082E-8
+ vbm = -3 dvtp0 = 0 dvtp1 = 0
+ dvt0 = 0 dvt1 = 0.53 dvt2 = -0.032
+ dvt0w = -3.58 dvt1w = 1.6706E6 dvt2w = 0.068
+ vfbsdoff = 0 u0 = 0.034334005492054 lu0 = -8.473052828464605E-9
+ wu0 = -2.144533275573204E-9 pu0 = 2.449109082616614E-15 ua = -1.319285758669252E-9
+ lua = 3.518420051115836E-15 wua = 3.107389201152689E-16 pua = -1.49618958209777E-21
+ ub = 3.129412952981256E-18 lub = -6.728708740039642E-24 wub = -7.36460815504153E-25
+ pub = 2.649401760059569E-30 uc = 1.534574804801472E-10 luc = -1.723693441454399E-16
+ wuc = -5.968161820187583E-17 puc = 1.024895154883428E-22 ud = 0
+ up = 0 lp = 1 eu = 1.67
+ vsat = 2.744759216612921E5 lvsat = -0.773262713250643 wvsat = -0.098459658570522
+ pvsat = 3.914889929899623E-7 a0 = 3.8297015144575 la0 = -9.646236747188062E-6
+ wa0 = -1.123489232311177E-6 pa0 = 4.117543055682662E-12 ags = 5.80339928648177E-3
+ lags = 2.120197132714229E-6 wags = 1.625088476121522E-7 pags = -9.236837358133756E-13
+ b0 = -7.069594045067998E-8 lb0 = 7.484216894700477E-13 wb0 = 3.61186422231201E-14
+ pb0 = -3.133978775515042E-19 b1 = -1.502706805526603E-8 lb1 = 4.497232457547178E-14
+ wb1 = 6.94655479516131E-15 pb1 = -1.340792229079888E-20 keta = 0.039148358622733
+ lketa = -1.41255661947602E-7 wketa = -1.95578945115152E-8 pketa = 7.601974717654816E-14
+ a1 = 0 a2 = 0.42385546 rdsw = 65.968
+ rdswmin = 0 rdw = 0 rdwmin = 0
+ rsw = 0 rswmin = 0 prwb = 0
+ prwg = 0.021507 wr = 1 voff = -0.211489952214131
+ lvoff = 2.749859149819424E-7 wvoff = 3.759180083987658E-8 pvoff = -1.012813113696829E-13
+ voffl = 5.8197729E-9 minv = 0 nfactor = 1.793296108457332
+ lnfactor = 2.96576296305798E-6 wnfactor = 3.785290273939828E-7 pnfactor = -7.97833841825676E-13
+ eta0 = 0.385916637942246 leta0 = -1.21636615712113E-6 weta0 = -1.151109243581842E-7
+ peta0 = 4.57696690333853E-13 etab = -0.337436557697938 letab = 1.06336412477885E-6
+ wetab = 1.006315628036956E-7 petab = -4.00124779600035E-13 dsub = 1.71440240732923
+ ldsub = -4.590060970268415E-6 wdsub = -4.343808466346573E-7 pdsub = 1.72715732201454E-12
+ cit = 0 cdsc = 0 cdscb = 0
+ cdscd = 5.4E-3 pclm = 6.524816574522276 lpclm = -1.928342377118752E-5
+ wpclm = -2.738217006099484E-6 ppclm = 9.15186121789064E-12 pdiblc1 = 0.39
+ pdiblc2 = 0.011484178912991 lpdiblc2 = -4.4170122448671E-8 wpdiblc2 = -4.561596409594461E-9
+ ppdiblc2 = 2.707069355309027E-14 pdiblcb = -0.073100100305385 lpdiblcb = 1.912525404278507E-7
+ wpdiblcb = 1.809920194311072E-8 ppdiblcb = -7.19648884172725E-14 drout = 0.56
+ pscbe1 = 1.124901769919126E8 lpscbe1 = 1.35861291159991E3 wpscbe1 = 258.6975712211291
+ ppscbe1 = -5.112215836026372E-4 pscbe2 = 1E-12 pvag = 0
+ delta = 0.01 fprout = 0 pdits = 0
+ pditsl = 0 pditsd = 0 lambda = 0
+ vtl = 0 lc = 5E-9 xn = 3
+ alpha0 = 3E-8 alpha1 = 0.85 beta0 = 13.86
+ aigbacc = 1 bigbacc = 0 cigbacc = 0
+ nigbacc = 0 aigbinv = 0.35 bigbinv = 0.03
+ cigbinv = 6E-3 eigbinv = 1.1 nigbinv = 0
+ aigc = 0.43 bigc = 0.054 cigc = 0.075
+ aigsd = 0.43 bigsd = 0.054 cigsd = 0.075
+ dlcig = 0 nigc = 0 poxedge = 1
+ pigcd = 1 ntox = 1 toxref = 4.148E-9
+ agidl = 0 bgidl = 2.3E9 cgidl = 0.5
+ egidl = 0.8 noia = 2.5E42 noib = 0
+ noic = 0 em = 4.1E7 af = 1
+ ef = 0.84 kf = 0 lintnoi = -1E-7
+ tnoia = 1.5E7 tnoib = 9.9E6 ntnoi = 1
+ rnoia = 0.94 rnoib = 0.26 xpart = 0
+ cgso = {2.449068E-10/sw_func_tox_lv_ratio} cgdo = {2.449068E-10/sw_func_tox_lv_ratio} cgbo = {1E-13/sw_func_tox_lv_ratio}
+ ckappas = 0.6 cf = 1.4067E-12 clc = 1E-7
+ cle = 0.6 dlc = 9.87908E-9 dwc = 0
+ vfbcv = -1 noff = 3.4037 voffcv = -0.17287
+ acde = 0.4 moin = 6.9 cgsl = {0/sw_func_tox_lv_ratio}
+ cgdl = {0/sw_func_tox_lv_ratio} ijthsrev = 0.1 ijthsfwd = 0.1
+ xjbvs = 1 bvs = 11.7 jss = 2.75E-3
+ jsws = 6E-10 cjs = {sw_nsd_pw_cj} mjs = 0.44
+ mjsws = 9E-4 cjsws = {3.67354204E-11*sw_func_nsd_pw_cj} cjswgs = {2.38232788E-10*sw_func_nsd_pw_cj}
+ mjswgs = 0.8 pbs = 0.729 pbsws = 0.2
+ pbswgs = 0.95578 xrcrg1 = 12 xrcrg2 = 1
+ rbpb = 50 rbpd = 50 rbps = 50
+ rbdb = 50 rbsb = 50 gbmin = 1E-12
+ tnom = 30 ute = 1.266885813638198 lute = -9.043810953278586E-6
+ wute = -1.083660424691519E-6 pute = 3.721448309833992E-12 kt1 = -0.122736454283736
+ lkt1 = -4.846815770746093E-7 wkt1 = -6.884135912113222E-8 pkt1 = 1.702401400398997E-13
+ kt1l = 0 kt2 = 0.10691246999792 lkt2 = -4.085959146185201E-7
+ wkt2 = -6.160097866040711E-8 pkt2 = 1.733447686553227E-13 ua1 = 9.276899010117521E-9
+ lua1 = -2.807868902479033E-14 wua1 = -3.613114343086065E-15 pua1 = 1.191767338145399E-20
+ ub1 = -5.964682768424203E-18 lub1 = 1.805071705310189E-23 wub1 = 2.267423394180929E-24
+ pub1 = -7.500929105687678E-30 uc1 = -1.35474356923058E-10 luc1 = 4.444956958484668E-16
+ wuc1 = 7.284972508210646E-17 puc1 = -1.768514161662088E-22 at = 2.578644857883144E5
+ lat = -0.468645225064405 wat = -0.044350284441399 pat = 1.763427625776845E-7
+ prt = 0 njs = 1.2928 xtis = 2
+ tpb = 1.2287E-3 tpbsw = 0 tpbswg = 0
+ tcj = 7.92E-4 tcjsw = 1E-5 tcjswg = 0
+ tvoff = 0 tvfbsdoff = 0 saref = 3E-6
+ sbref = 3E-6 wlod = 0 ku0 = -2.7E-8
+ kvsat = 0.2 kvth0 = 9.8E-9 tku0 = 0
+ llodku0 = 0 wlodku0 = 1 llodvth = 0
+ wlodvth = 1 lku0 = 0 wku0 = 0
+ pku0 = 0 lkvth0 = 0 wkvth0 = 2E-7
+ pkvth0 = 0 stk2 = 0 lodk2 = 1
+ steta0 = 0 lodeta0 = 1

.model nshort_model.44 nmos
+ level = 54 lmin = 1E-6 lmax = 2E-6 wmin = 4.2E-7
+ wmax = 5.5E-7 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 4.148E-9
+ toxm = 4.148E-9 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 9.999999999999999E22 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {2.1859E-8+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {1.1932E-8-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = 0 dwb = 0 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = 0.458352341089585 lvth0 = 1.608157758219257E-7
+ wvth0 = 1.335813477926378E-8 pvth0 = -4.786007491003511E-14 k1 = 0.504278926725039
+ lk1 = -4.009620621353525E-8 wk1 = 4.418761684959186E-8 pk1 = 1.832337479412715E-15
+ k2 = -9.235621793401759E-3 lk2 = 1.414505904470154E-8 wk2 = -2.063800994412376E-8
+ pk2 = -2.053172858231422E-15 k3 = 2 k3b = 0.54
+ w0 = 0 lpe0 = 1.0325E-7 lpeb = -7.082E-8
+ vbm = -3 dvtp0 = 0 dvtp1 = 0
+ dvt0 = 0 dvt1 = 0.53 dvt2 = -0.032
+ dvt0w = -3.58 dvt1w = 1.6706E6 dvt2w = 0.068
+ vfbsdoff = 0 u0 = 0.028240903287362 lu0 = 3.56774578990764E-9
+ wu0 = 1.324023540467803E-9 pu0 = -4.405230909607398E-15 ua = 1.759826551584098E-9
+ lua = -2.566324633218979E-15 wua = -7.515159048925582E-16 pua = 6.029704187738978E-22
+ ub = -2.469591411946504E-18 lub = 4.33568534965124E-24 wub = 1.2814326832801E-24
+ pub = -1.33823022705395E-30 uc = 1.007167048325207E-10 luc = -6.814639872024185E-17
+ wuc = -1.972366560568082E-17 puc = 2.352716687670837E-23 ud = 0
+ up = 0 lp = 1 eu = 1.67
+ vsat = -5.069920090094171E4 lvsat = -0.130672447251001 wvsat = 0.064482465335552
+ pvsat = 6.949319602270801E-8 a0 = -2.401967977478693 la0 = 2.668389675928758E-6
+ wa0 = 1.468240314501637E-6 pa0 = -1.004067004037825E-12 ags = -2.048764178011694
+ lags = 6.180302086645936E-6 wags = 8.96182007674527E-7 pags = -2.373521679646397E-12
+ b0 = -4.790817907314026E-7 lb0 = 1.555447670100394E-12 wb0 = 2.522826007216898E-13
+ pb0 = -7.405672578430336E-19 b1 = 2.089263969396732E-8 lb1 = -2.600990301726723E-14
+ wb1 = -3.612608292866927E-15 pb1 = 7.458420017324892E-21 keta = 0.224654549095109
+ lketa = -5.078411231629214E-7 wketa = -7.774035724088573E-8 pketa = 1.909962063447155E-13
+ a1 = 0 a2 = 0.42385546 rdsw = 65.968
+ rdswmin = 0 rdw = 0 rdwmin = 0
+ rsw = 0 rswmin = 0 prwb = 0
+ prwg = 0.021507 wr = 1 voff = 0.031168115482247
+ lvoff = -2.045394282833073E-7 wvoff = -4.8594048803842E-8 pvoff = 6.903364880185656E-14
+ voffl = 5.8197729E-9 minv = 0 nfactor = 4.865453049045523
+ lnfactor = -3.105236964888206E-6 wnfactor = -6.410805266612126E-7 pnfactor = 1.217053303886742E-12
+ eta0 = -0.456213240134492 leta0 = 4.477970116219225E-7 weta0 = 2.302218487163684E-7
+ peta0 = -2.24727834518601E-13 etab = 0.716415520657146 letab = -1.019190905933453E-6
+ wetab = -3.215103913865672E-7 petab = 4.34085133185694E-13 dsub = -1.455964014658461
+ ldsub = 1.675014249412651E-6 wdsub = 8.687616932693149E-7 pdsub = -8.48029564221136E-13
+ cit = 0 cdsc = 0 cdscb = 0
+ cdscd = 5.4E-3 pclm = -6.772708011175367 lpclm = 6.994293273494672E-6
+ wpclm = 3.504661816301313E-6 ppclm = -3.184916366693179E-12 pdiblc1 = 1.088856024828547
+ lpdiblc1 = -1.381034549480586E-6 wpdiblc1 = -3.362090663973831E-7 ppdiblc1 = 6.643948396342592E-13
+ pdiblc2 = -0.022827071647606 lpdiblc2 = 2.363357498914499E-8 wpdiblc2 = 1.642038104829278E-8
+ ppdiblc2 = -1.439254745262919E-14 pdiblcb = -0.023110275910473 lpdiblcb = 9.246584880738681E-8
+ wpdiblcb = -7.110691598555593E-10 ppdiblcb = -3.479323452094112E-14 drout = -0.541207011951394
+ ldrout = 2.17613481976958E-6 wdrout = 3.797557777796574E-7 pdrout = -7.504490636783811E-13
+ pscbe1 = 1.051292570600871E9 lpscbe1 = -496.5882952969237 wpscbe1 = -94.55687105083712
+ ppscbe1 = 1.86857236930917E-4 pscbe2 = 1E-12 pvag = 0
+ delta = 0.01 fprout = 0 pdits = 0
+ pditsl = 0 pditsd = 0 lambda = 0
+ vtl = 0 lc = 5E-9 xn = 3
+ alpha0 = -2.084044980055752E-5 lalpha0 = 4.124284718707455E-11 walpha0 = 7.853174591853387E-12
+ palpha0 = -1.551894102524679E-17 alpha1 = 0.85 beta0 = 0.159252990672252
+ lbeta0 = 2.70745393920249E-5 wbeta0 = 5.155344486163863E-6 pbeta0 = -1.018766183150991E-11
+ aigbacc = 1 bigbacc = 0 cigbacc = 0
+ nigbacc = 0 aigbinv = 0.35 bigbinv = 0.03
+ cigbinv = 6E-3 eigbinv = 1.1 nigbinv = 0
+ aigc = 0.43 bigc = 0.054 cigc = 0.075
+ aigsd = 0.43 bigsd = 0.054 cigsd = 0.075
+ dlcig = 0 nigc = 0 poxedge = 1
+ pigcd = 1 ntox = 1 toxref = 4.148E-9
+ agidl = 0 bgidl = 2.3E9 cgidl = 0.5
+ egidl = 0.8 noia = 2.5E42 noib = 0
+ noic = 0 em = 4.1E7 af = 1
+ ef = 0.84 kf = 0 lintnoi = -1E-7
+ tnoia = 1.5E7 tnoib = 9.9E6 ntnoi = 1
+ rnoia = 0.94 rnoib = 0.26 xpart = 0
+ cgso = {2.449068E-10/sw_func_tox_lv_ratio} cgdo = {2.449068E-10/sw_func_tox_lv_ratio} cgbo = {1E-13/sw_func_tox_lv_ratio}
+ ckappas = 0.6 cf = 1.4067E-12 clc = 1E-7
+ cle = 0.6 dlc = 9.87908E-9 dwc = 0
+ vfbcv = -1 noff = 3.4037 voffcv = -0.17287
+ acde = 0.4 moin = 6.9 cgsl = {0/sw_func_tox_lv_ratio}
+ cgdl = {0/sw_func_tox_lv_ratio} ijthsrev = 0.1 ijthsfwd = 0.1
+ xjbvs = 1 bvs = 11.7 jss = 2.75E-3
+ jsws = 6E-10 cjs = {sw_nsd_pw_cj} mjs = 0.44
+ mjsws = 9E-4 cjsws = {3.67354204E-11*sw_func_nsd_pw_cj} cjswgs = {2.38232788E-10*sw_func_nsd_pw_cj}
+ mjswgs = 0.8 pbs = 0.729 pbsws = 0.2
+ pbswgs = 0.95578 xrcrg1 = 12 xrcrg2 = 1
+ rbpb = 50 rbpd = 50 rbps = 50
+ rbdb = 50 rbsb = 50 gbmin = 1E-12
+ tnom = 30 ute = -4.486928109870582 lute = 2.326507878268359E-6
+ wute = 1.071488941632694E-6 pute = -5.374199383364716E-13 kt1 = -0.519358627898
+ lkt1 = 2.990977786027869E-7 wkt1 = 6.469651778461342E-8 pkt1 = -9.364886587711284E-14
+ kt1l = 0 kt2 = -0.168959029967806 lkt2 = 1.365636878377489E-7
+ wkt2 = 5.065862628426374E-8 pkt2 = -4.849547802161935E-14 ua1 = -8.418260372782712E-9
+ lua1 = 6.889352457496604E-15 wua1 = 3.471969351903148E-15 pua1 = -2.083415571227209E-21
+ ub1 = 4.961522835964977E-18 lub1 = -3.540951185133325E-24 wub1 = -2.029634320913872E-24
+ pub1 = 9.906413391889016E-31 uc1 = 1.55239391369662E-10 luc1 = -1.299942078477158E-16
+ wuc1 = -4.225474315696772E-17 puc1 = 5.061066728188228E-23 at = 1.699214760120113E5
+ lat = -0.294857877497101 wat = -7.585888773231654E-3 pat = 1.036913167795759E-7
+ prt = 0 njs = 1.2928 xtis = 2
+ tpb = 1.2287E-3 tpbsw = 0 tpbswg = 0
+ tcj = 7.92E-4 tcjsw = 1E-5 tcjswg = 0
+ tvoff = 0 tvfbsdoff = 0 saref = 3E-6
+ sbref = 3E-6 wlod = 0 ku0 = -2.7E-8
+ kvsat = 0.2 kvth0 = 9.8E-9 tku0 = 0
+ llodku0 = 0 wlodku0 = 1 llodvth = 0
+ wlodvth = 1 lku0 = 0 wku0 = 0
+ pku0 = 0 lkvth0 = 0 wkvth0 = 2E-7
+ pkvth0 = 0 stk2 = 0 lodk2 = 1
+ steta0 = 0 lodeta0 = 1

.model nshort_model.45 nmos
+ level = 54 lmin = 5E-7 lmax = 1E-6 wmin = 4.2E-7
+ wmax = 5.5E-7 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 4.148E-9
+ toxm = 4.148E-9 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 9.999999999999999E22 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {2.1859E-8+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {1.1932E-8-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = 0 dwb = 0 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = 0.602075679641821 lvth0 = 2.052225102090036E-8
+ wvth0 = -3.245887471432459E-8 pvth0 = -3.136442531001726E-15 k1 = 0.729032643201111
+ lk1 = -2.59486399999622E-7 wk1 = -5.033422151606413E-8 pk1 = 9.409850669431069E-14
+ k2 = -0.081367191490095 lk2 = 8.455528096215271E-8 wk2 = 6.589730746570213E-9
+ pk2 = -2.863115074508267E-14 k3 = 2 k3b = 0.54
+ w0 = 0 lpe0 = 1.0325E-7 lpeb = -7.082E-8
+ vbm = -3 dvtp0 = 0 dvtp1 = 0
+ dvt0 = 0 dvt1 = 0.53 dvt2 = -0.032
+ dvt0w = -3.58 dvt1w = 1.6706E6 dvt2w = 0.068
+ vfbsdoff = 0 u0 = 0.047557179028213 lu0 = -1.528756634666354E-8
+ wu0 = -9.11218586846113E-9 pu0 = 5.781928797986857E-15 ua = 4.871857930411846E-10
+ lua = -1.324054173737934E-15 wua = -6.670888867208654E-16 pua = 5.205581669638543E-22
+ ub = 1.159843505751688E-18 lub = 7.928632668289976E-25 wub = 2.729428420073434E-25
+ pub = -3.538069873533256E-31 uc = -1.223667895511096E-10 luc = 1.496134311534176E-16
+ wuc = 7.571725253912618E-17 puc = -6.963614919749097E-23 ud = 0
+ up = 0 lp = 1 eu = 1.67
+ vsat = -5.043837954004782E5 lvsat = 0.312185418085398 wvsat = 0.254921140785259
+ pvsat = -1.164008508760673E-7 a0 = -0.352950882162756 la0 = 6.682703245754402E-7
+ wa0 = 6.972320638419662E-7 pa0 = -2.514580942718958E-13 ags = 7.835224833576818
+ lags = -3.467815411170028E-6 wags = -2.806664047797939E-6 pags = 1.240959657558274E-12
+ b0 = 2.17559737444601E-6 lb0 = -1.035880231479226E-12 wb0 = -9.886102582099323E-13
+ pb0 = 4.707129339030443E-19 b1 = -1.123169055391349E-8 lb1 = 5.347812213578154E-15
+ wb1 = 7.864046017517882E-15 pb1 = -3.744355414596895E-21 keta = -0.555539398388321
+ lketa = 2.53734275957764E-7 wketa = 2.227381012765366E-7 pketa = -1.02311634238647E-13
+ a1 = 0 a2 = 0.42385546 rdsw = 65.968
+ rdswmin = 0 rdw = 0 rdwmin = 0
+ rsw = 0 rswmin = 0 prwb = 0
+ prwg = 0.021507 wr = 1 voff = -0.18244212567183
+ lvoff = 3.973218075868783E-9 wvoff = 2.851270325730272E-8 pvoff = -6.233027728101018E-15
+ voffl = 5.8197729E-9 minv = 0 nfactor = 1.869806735684398
+ lnfactor = -1.810787551491305E-7 wnfactor = 4.623731158037607E-7 pnfactor = 1.399324791455524E-13
+ eta0 = -0.4616715915 leta0 = 4.531251048904439E-7 etab = -0.638287327607384
+ letab = 3.031833135600926E-7 wetab = 2.400584440817618E-7 petab = -1.140824235930188E-13
+ dsub = 0.198081081154105 ldsub = 6.044128576655695E-8 wdsub = 7.094452481555044E-9
+ pdsub = -6.925150467535216E-15 cit = 0 cdsc = 0
+ cdscb = 0 cdscd = 5.4E-3 pclm = 0.802973974241045
+ lpclm = -4.00602637021765E-7 wpclm = 2.358871250751005E-7 ppclm = 5.852285301611672E-15
+ pdiblc1 = 0.618462828466831 lpdiblc1 = -9.218668163568458E-7 wpdiblc1 = 2.12159228206922E-8
+ ppdiblc1 = 3.154994403588839E-13 pdiblc2 = 6.182493560126774E-3 lpdiblc2 = -4.68370595447023E-9
+ wpdiblc2 = 1.487707263858081E-9 ppdiblc2 = 1.837730046137614E-16 pdiblcb = 0.421758927318469
+ lpdiblcb = -3.417869957556997E-7 wpdiblcb = -1.681073426892483E-7 ppdiblcb = 1.286082943369462E-13
+ drout = 2.343414714762921 ldrout = -6.396482940584242E-7 wdrout = -7.595116951073072E-7
+ pdrout = 3.61630930235609E-13 pscbe1 = 1.643833659825361E9 lpscbe1 = -1.07498898396816E3
+ wpscbe1 = -317.5194171864063 ppscbe1 = 4.04499004865507E-4 pscbe2 = 1E-12
+ pvag = 0 delta = 0.01 fprout = 0
+ pdits = 0 pditsl = 0 pditsd = 0
+ lambda = 0 vtl = 0 lc = 5E-9
+ xn = 3 alpha0 = 2.898972017709044E-5 lalpha0 = -7.39817561422683E-12
+ walpha0 = -1.110126543091722E-11 palpha0 = 2.98317024082043E-18 alpha1 = 0.85
+ beta0 = 30.637142726361084 lbeta0 = -2.676025983011462E-6 wbeta0 = -6.936418513465561E-6
+ pbeta0 = 1.615543335896358E-12 aigbacc = 1 bigbacc = 0
+ cigbacc = 0 nigbacc = 0 aigbinv = 0.35
+ bigbinv = 0.03 cigbinv = 6E-3 eigbinv = 1.1
+ nigbinv = 0 aigc = 0.43 bigc = 0.054
+ cigc = 0.075 aigsd = 0.43 bigsd = 0.054
+ cigsd = 0.075 dlcig = 0 nigc = 0
+ poxedge = 1 pigcd = 1 ntox = 1
+ toxref = 4.148E-9 agidl = 0 bgidl = 2.3E9
+ cgidl = 0.5 egidl = 0.8 noia = 2.5E42
+ noib = 0 noic = 0 em = 4.1E7
+ af = 1 ef = 0.84 kf = 0
+ lintnoi = -1E-7 tnoia = 1.5E7 tnoib = 9.9E6
+ ntnoi = 1 rnoia = 0.94 rnoib = 0.26
+ xpart = 0 cgso = {2.449068E-10/sw_func_tox_lv_ratio} cgdo = {2.449068E-10/sw_func_tox_lv_ratio}
+ cgbo = {1E-13/sw_func_tox_lv_ratio} ckappas = 0.6 cf = 1.4067E-12
+ clc = 1E-7 cle = 0.6 dlc = 9.87908E-9
+ dwc = 0 vfbcv = -1 noff = 3.4037
+ voffcv = -0.17287 acde = 0.4 moin = 6.9
+ cgsl = {0/sw_func_tox_lv_ratio} cgdl = {0/sw_func_tox_lv_ratio} ijthsrev = 0.1
+ ijthsfwd = 0.1 xjbvs = 1 bvs = 11.7
+ jss = 2.75E-3 jsws = 6E-10 cjs = {sw_nsd_pw_cj}
+ mjs = 0.44 mjsws = 9E-4 cjsws = {3.67354204E-11*sw_func_nsd_pw_cj}
+ cjswgs = {2.38232788E-10*sw_func_nsd_pw_cj} mjswgs = 0.8 pbs = 0.729
+ pbsws = 0.2 pbswgs = 0.95578 xrcrg1 = 12
+ xrcrg2 = 1 rbpb = 50 rbpd = 50
+ rbps = 50 rbdb = 50 rbsb = 50
+ gbmin = 1E-12 tnom = 30 ute = -3.339164895010054
+ lute = 1.206134884767262E-6 wute = 1.260123937306694E-6 pute = -7.21553348473707E-13
+ kt1 = -0.224164772045984 lkt1 = 1.094842892682366E-8 wkt1 = -2.349379509523284E-8
+ pkt1 = -7.563126623831228E-15 kt1l = 0 kt2 = -0.058042814665814
+ lkt2 = 2.829437709772421E-8 wkt2 = 2.02775378525433E-8 pkt2 = -1.883940388423349E-14
+ ua1 = -4.6966301439315E-9 lua1 = 3.256535212426696E-15 wua1 = 3.243553972719166E-15
+ pua1 = -1.860451096652075E-21 ub1 = 5.09380394287127E-18 lub1 = -3.670075535704408E-24
+ wub1 = -2.936846143416803E-24 pub1 = 1.876203458759623E-30 uc1 = 3.148457653824608E-10
+ luc1 = -2.85791735351073E-16 wuc1 = -1.216285396991255E-16 puc1 = 1.28090287543358E-22
+ at = -2.974989265687112E5 lat = 0.161408004596435 wat = 0.207442116738648
+ pat = -1.06205260408768E-7 prt = 0 njs = 1.2928
+ xtis = 2 tpb = 1.2287E-3 tpbsw = 0
+ tpbswg = 0 tcj = 7.92E-4 tcjsw = 1E-5
+ tcjswg = 0 tvoff = 0 tvfbsdoff = 0
+ saref = 2.75E-6 sbref = 2.74E-6 wlod = 0
+ ku0 = -2.7E-8 kvsat = 0.2 kvth0 = 9.8E-9
+ tku0 = 0 llodku0 = 0 wlodku0 = 1
+ llodvth = 0 wlodvth = 1 lku0 = 0
+ wku0 = 0 pku0 = 0 lkvth0 = 0
+ wkvth0 = 2E-7 pkvth0 = 0 stk2 = 0
+ lodk2 = 1 steta0 = 0 lodeta0 = 1

.model nshort_model.46 nmos
+ level = 54 lmin = 2.5E-7 lmax = 5E-7 wmin = 4.2E-7
+ wmax = 5.5E-7 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 4.148E-9
+ toxm = 4.148E-9 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 9.999999999999999E22 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {2.1859E-8+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {1.1932E-8-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = 0 dwb = 0 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = 0.67972630614978 lvth0 = -1.645000768209284E-8
+ wvth0 = -3.361654371616982E-8 pvth0 = -2.585234643139145E-15 k1 = -0.076520957517309
+ lk1 = 1.240666692320434E-7 wk1 = 2.003787765672515E-7 pk1 = -2.527497736108685E-14
+ k2 = 0.173761406632363 lk2 = -3.692062923348205E-8 wk2 = -7.024308344881233E-8
+ pk2 = 7.951718074649985E-15 k3 = 2 k3b = 0.54
+ w0 = 0 lpe0 = 1.0325E-7 lpeb = -7.082E-8
+ vbm = -3 dvtp0 = 0 dvtp1 = 0
+ dvt0 = 0 dvt1 = 0.53 dvt2 = -0.032
+ dvt0w = -3.58 dvt1w = 1.6706E6 dvt2w = 0.068
+ vfbsdoff = 0 u0 = 0.018026142414072 lu0 = -1.226776697352957E-9
+ wu0 = 9.875938313578809E-10 pu0 = 9.730600908338322E-16 ua = -2.720006857721899E-9
+ lua = 2.030057062257979E-16 wua = 5.917959814325434E-16 pua = -7.884223861923712E-23
+ ub = 3.535966276517203E-18 lub = -3.384943247522118E-25 wub = -8.950130789557861E-25
+ pub = 2.022988730303751E-31 uc = 2.093837036698901E-10 luc = -8.344921686856368E-18
+ wuc = -8.57886803404576E-17 puc = 7.262639660062531E-24 ud = 0
+ up = 0 lp = 1 eu = 1.67
+ vsat = 1.488410930614433E5 lvsat = 1.161532592693065E-3 wvsat = 9.435089738563654E-3
+ pvsat = 4.838955251021425E-10 a0 = 0.888610580988555 la0 = 7.711821575642732E-8
+ wa0 = 2.300548333644644E-7 pa0 = -2.901819646125998E-14 ags = 0.300420571971155
+ lags = 1.197761507338455E-7 wags = -2.725546728687004E-7 pags = 3.437895621696669E-14
+ b0 = 0 b1 = 0 keta = -0.089285003730642
+ lketa = 3.17337735030355E-8 wketa = 4.523053790070627E-8 pketa = -1.77938930431327E-14
+ a1 = 0 a2 = 0.42385546 rdsw = 65.968
+ rdswmin = 0 rdw = 0 rdwmin = 0
+ rsw = 0 rswmin = 0 prwb = 0
+ prwg = 0.021507 wr = 1 voff = -0.162048690837183
+ lvoff = -5.736830412560864E-9 wvoff = 2.097970500005218E-8 pvoff = -2.646296069886775E-15
+ voffl = 5.8197729E-9 minv = 0 nfactor = 0.748455796562336
+ lnfactor = 3.528367956006915E-7 wnfactor = 1.192177911767006E-6 pnfactor = -2.075538571852033E-13
+ eta0 = 0.665616158886314 leta0 = -8.36171754274942E-8 weta0 = 3.665893947397869E-10
+ peta0 = -1.745464080538232E-16 etab = 0.013775629344064 letab = -7.287334510942259E-9
+ wetab = 6.22982109414962E-10 petab = -7.858047135344273E-17 dsub = 0.449100370013342
+ ldsub = -5.907803435372468E-8 wdsub = -9.733034860537417E-8 pdsub = 4.27952566227909E-14
+ cit = 0 cdsc = 0 cdscb = 0
+ cdscd = 6.606580937142858E-3 lcdscd = -5.744966210874517E-10 pclm = -0.131544499626994
+ lpclm = 4.43552510518678E-8 wpclm = 3.479701394640708E-7 ppclm = -4.751447283749513E-14
+ pdiblc1 = -1.921204109069609 lpdiblc1 = 2.873600406140047E-7 wpdiblc1 = 9.302888713915348E-7
+ ppdiblc1 = -1.173429170818428E-13 pdiblc2 = -8.000890161632314E-3 lpdiblc2 = 2.069513637273254E-9
+ wpdiblc2 = 2.548925686851695E-9 ppdiblc2 = -3.215112904367258E-16 pdiblcb = -0.365551633980779
+ lpdiblcb = 3.307990565907937E-8 wpdiblcb = 1.387609617664519E-7 ppdiblcb = -1.750275267337307E-14
+ drout = 1.178994865669069 ldrout = -8.52260847902744E-8 pdrout = -1.110048380034836E-19
+ pscbe1 = -1.120363252849234E9 lpscbe1 = 241.14467724507114 wpscbe1 = 723.7616561258297
+ ppscbe1 = -9.129240025708776E-5 pscbe2 = 1E-12 pvag = 0
+ delta = 0.01 fprout = 0 pdits = 0
+ pditsl = 0 pditsd = 0 lambda = 0
+ vtl = 0 lc = 5E-9 xn = 3
+ alpha0 = 1.82888277486066E-5 lalpha0 = -2.303095496898244E-12 walpha0 = -6.578691075413642E-12
+ palpha0 = 8.298097774883765E-19 alpha1 = 0.85 beta0 = 29.041248588991984
+ lbeta0 = -1.916163332021091E-6 wbeta0 = -4.820386369803083E-6 pbeta0 = 6.080242551414806E-13
+ aigbacc = 1 bigbacc = 0 cigbacc = 0
+ nigbacc = 0 aigbinv = 0.35 bigbinv = 0.03
+ cigbinv = 6E-3 eigbinv = 1.1 nigbinv = 0
+ aigc = 0.43 bigc = 0.054 cigc = 0.075
+ aigsd = 0.43 bigsd = 0.054 cigsd = 0.075
+ dlcig = 0 nigc = 0 poxedge = 1
+ pigcd = 1 ntox = 1 toxref = 4.148E-9
+ agidl = 0 bgidl = 2.3E9 cgidl = 0.5
+ egidl = 0.8 noia = 2.5E42 noib = 0
+ noic = 0 em = 4.1E7 af = 1
+ ef = 0.84 kf = 0 lintnoi = -1E-7
+ tnoia = 1.5E7 tnoib = 9.9E6 ntnoi = 1
+ rnoia = 0.94 rnoib = 0.26 xpart = 0
+ cgso = {2.449068E-10/sw_func_tox_lv_ratio} cgdo = {2.449068E-10/sw_func_tox_lv_ratio} cgbo = {1E-13/sw_func_tox_lv_ratio}
+ ckappas = 0.6 cf = 1.4067E-12 clc = 1E-7
+ cle = 0.6 dlc = 9.87908E-9 dwc = 0
+ vfbcv = -1 noff = 3.4037 voffcv = -0.17287
+ acde = 0.4 moin = 6.9 cgsl = {0/sw_func_tox_lv_ratio}
+ cgdl = {0/sw_func_tox_lv_ratio} ijthsrev = 0.1 ijthsfwd = 0.1
+ xjbvs = 1 bvs = 11.7 jss = 2.75E-3
+ jsws = 6E-10 cjs = {sw_nsd_pw_cj} mjs = 0.44
+ mjsws = 9E-4 cjsws = {3.67354204E-11*sw_func_nsd_pw_cj} cjswgs = {2.38232788E-10*sw_func_nsd_pw_cj}
+ mjswgs = 0.8 pbs = 0.729 pbsws = 0.2
+ pbswgs = 0.95578 xrcrg1 = 12 xrcrg2 = 1
+ rbpb = 50 rbpd = 50 rbps = 50
+ rbdb = 50 rbsb = 50 gbmin = 1E-12
+ tnom = 30 ute = -0.60660595407415 lute = -9.493479913419512E-8
+ wute = -3.663351553875833E-7 pute = 5.286237808537516E-14 kt1 = -0.186830471644066
+ lkt1 = -6.827775529343827E-9 wkt1 = -5.356962355798546E-8 pkt1 = 6.757058037109957E-15
+ kt1l = 0 kt2 = 0.012287935267732 lkt2 = -5.192624852634505E-9
+ wkt2 = -2.624153748935701E-8 pkt2 = 3.310002572757552E-15 ua1 = 2.923738656541207E-9
+ lua1 = -3.717967067551776E-16 wua1 = -9.030808065641764E-16 pua1 = 1.139110006167789E-22
+ ub1 = -3.811443586893063E-18 lub1 = 5.700334021274635E-25 wub1 = 1.365329381193485E-24
+ pub1 = -1.722171868262214E-31 uc1 = -4.412794766712278E-10 luc1 = 7.422671289940197E-17
+ wuc1 = 2.005101747576434E-16 puc1 = -2.529155140323011E-23 at = 3.709133813566698E4
+ lat = 2.097534321151525E-3 wat = -0.0212417163237 pat = 2.67934513020611E-9
+ prt = 0 njs = 1.2928 xtis = 2
+ tpb = 1.2287E-3 tpbsw = 0 tpbswg = 0
+ tcj = 7.92E-4 tcjsw = 1E-5 tcjswg = 0
+ tvoff = 0 tvfbsdoff = 0 saref = 1.75E-6
+ sbref = 1.74E-6 wlod = 0 ku0 = -2.7E-8
+ kvsat = 0.2 kvth0 = 9.8E-9 tku0 = 0
+ llodku0 = 0 wlodku0 = 1 llodvth = 0
+ wlodvth = 1 lku0 = 0 wku0 = 0
+ pku0 = 0 lkvth0 = 0 wkvth0 = 2E-7
+ pkvth0 = 0 stk2 = 0 lodk2 = 1
+ steta0 = 0 lodeta0 = 1

.model nshort_model.47 nmos
+ level = 54 lmin = 1.8E-7 lmax = 2.5E-7 wmin = 4.2E-7
+ wmax = 5.5E-7 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 4.148E-9
+ toxm = 4.148E-9 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 9.999999999999999E22 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {2.1859E-8+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {1.1932E-8-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = 0 dwb = 0 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = 0.703442596798674 lvth0 = -2.181311478427132E-8
+ wvth0 = -4.562367477847243E-8 pvth0 = 1.300099467657357E-16 k1 = 0.483028853472105
+ lk1 = -2.467686825858748E-9 wk1 = -8.29112208400912E-8 pk1 = 3.878708949261999E-14
+ k2 = -0.016012976078611 lk2 = 5.99419057524682E-9 wk2 = 2.583627057886455E-8
+ pk2 = -1.377528272775275E-14 k3 = 2 k3b = 0.54
+ w0 = 0 lpe0 = 1.0325E-7 lpeb = -7.082E-8
+ vbm = -3 dvtp0 = 0 dvtp1 = 0
+ dvt0 = 0 dvt1 = 0.53 dvt2 = -0.032
+ dvt0w = -3.58 dvt1w = 1.6706E6 dvt2w = 0.068
+ vfbsdoff = 0 u0 = -0.014343464950447 lu0 = 6.093156833629849E-9
+ wu0 = 1.737574338708012E-8 pu0 = -2.732890497098971E-15 ua = -2.565002500934947E-9
+ lua = 1.679536409994237E-16 wua = 5.133200656697319E-16 pua = -6.109600893229798E-23
+ ub = 3.348181225607259E-19 lub = 3.854005141908902E-25 wub = 7.256706107256089E-25
+ pub = -1.641960538194169E-31 uc = 4.669542172334981E-10 luc = -6.659088734207638E-17
+ wuc = -2.161919950884681E-16 puc = 3.675152364391862E-23 ud = 0
+ up = 0 lp = 1 eu = 1.67
+ vsat = 1.113617015379312E5 lvsat = 9.636972274254006E-3 wvsat = 0.02841023103787
+ pvsat = -3.807067027757848E-9 a0 = 0.888610580988552 la0 = 7.711821575642798E-8
+ wa0 = 2.300548333644655E-7 pa0 = -2.901819646126023E-14 ags = 2.376896349574169
+ lags = -3.497897757101894E-7 wags = -1.32383698250511E-6 pags = 2.721117325889058E-13
+ b0 = 0 b1 = 0 keta = -0.087157710034774
+ lketa = 3.125271581582667E-8 wketa = 4.415352739377523E-8 pketa = -1.755034219513734E-14
+ a1 = 0 a2 = 0.42385546 rdsw = 65.968
+ rdswmin = 0 rdw = 0 rdwmin = 0
+ rsw = 0 rswmin = 0 prwb = 0
+ prwg = 0.021507 wr = 1 voff = -0.287631667676037
+ lvoff = 2.26620016378703E-8 wvoff = 8.456010567998105E-8 pvoff = -1.702411355804317E-14
+ voffl = 5.8197729E-9 minv = 0 nfactor = -9.458934841244606
+ lnfactor = 2.661095284871801E-6 wnfactor = 6.359996058657179E-6 pnfactor = -1.376183581650359E-12
+ eta0 = -0.161282639661378 leta0 = 1.033744112808867E-7 weta0 = 4.190105669210626E-7
+ peta0 = -9.484502090994637E-14 etab = -0.059945773643593 letab = 9.383728675074594E-9
+ wetab = 3.794680145681231E-8 petab = -8.518839683296487E-15 dsub = 0.986595980022171
+ ldsub = -1.806251416186813E-7 wdsub = -3.69454701031865E-7 pdsub = 1.043323691831078E-13
+ cit = 0 cdsc = 0 cdscb = 0
+ cdscd = 9.566683299231139E-4 lcdscd = 7.031520162587922E-10 wcdscd = 2.860449054608426E-9
+ pcdscd = -6.468505074129308E-16 pclm = -0.695842177563804 lpclm = 1.719632707497862E-7
+ wpclm = 6.33663896445275E-7 ppclm = -1.121201162661967E-13 pdiblc1 = -2.162035380310168
+ lpdiblc1 = 3.418206609672597E-7 wpdiblc1 = 1.052217409057748E-6 ppdiblc1 = -1.449153488755296E-13
+ pdiblc2 = 3.948782161971526E-3 lpdiblc2 = -6.327374632972238E-10 wpdiblc2 = -3.500978316487108E-9
+ ppdiblc2 = 1.046589801262298E-15 pdiblcb = -0.497679548561119 lpdiblcb = 6.295878375061909E-8
+ wpdiblcb = 2.056549466160158E-7 ppdiblcb = -3.262989083131406E-14 drout = 0.340837902238698
+ ldrout = 1.043113782920161E-7 wdrout = 4.243437837594535E-7 pdrout = -9.595943102997833E-14
+ pscbe1 = -1.134842622072485E9 lpscbe1 = 244.41898388374022 wpscbe1 = 731.0923001349155
+ ppscbe1 = -9.295012277072637E-5 pscbe2 = 1E-12 pvag = 0
+ delta = 0.01 fprout = 0 pdits = 0
+ pditsl = 0 pditsd = 0 lambda = 0
+ vtl = 0 lc = 5E-9 xn = 3
+ alpha0 = 1.746637838251613E-5 lalpha0 = -2.117110087048012E-12 walpha0 = -6.162299765450633E-12
+ palpha0 = 7.356487122185814E-19 alpha1 = 0.85 beta0 = 29.638933263805214
+ lbeta0 = -2.051321353644654E-6 wbeta0 = -5.122983362336866E-6 pbeta0 = 6.764523286451002E-13
+ aigbacc = 1 bigbacc = 0 cigbacc = 0
+ nigbacc = 0 aigbinv = 0.35 bigbinv = 0.03
+ cigbinv = 6E-3 eigbinv = 1.1 nigbinv = 0
+ aigc = 0.43 bigc = 0.054 cigc = 0.075
+ aigsd = 0.43 bigsd = 0.054 cigsd = 0.075
+ dlcig = 0 nigc = 0 poxedge = 1
+ pigcd = 1 ntox = 1 toxref = 4.148E-9
+ agidl = 0 bgidl = 2.3E9 cgidl = 0.5
+ egidl = 0.8 noia = 2.5E42 noib = 0
+ noic = 0 em = 4.1E7 af = 1
+ ef = 0.84 kf = 0 lintnoi = -1E-7
+ tnoia = 1.5E7 tnoib = 9.9E6 ntnoi = 1
+ rnoia = 0.94 rnoib = 0.26 xpart = 0
+ cgso = {2.449068E-10/sw_func_tox_lv_ratio} cgdo = {2.449068E-10/sw_func_tox_lv_ratio} cgbo = {1E-13/sw_func_tox_lv_ratio}
+ ckappas = 0.6 cf = 1.4067E-12 clc = 1E-7
+ cle = 0.6 dlc = 9.87908E-9 dwc = 0
+ vfbcv = -1 noff = 3.4037 voffcv = -0.17287
+ acde = 0.4 moin = 6.9 cgsl = {0/sw_func_tox_lv_ratio}
+ cgdl = {0/sw_func_tox_lv_ratio} ijthsrev = 0.1 ijthsfwd = 0.1
+ xjbvs = 1 bvs = 11.7 jss = 2.75E-3
+ jsws = 6E-10 cjs = {sw_nsd_pw_cj} mjs = 0.44
+ mjsws = 9E-4 cjsws = {3.67354204E-11*sw_func_nsd_pw_cj} cjswgs = {2.38232788E-10*sw_func_nsd_pw_cj}
+ mjswgs = 0.8 pbs = 0.729 pbsws = 0.2
+ pbswgs = 0.95578 xrcrg1 = 12 xrcrg2 = 1
+ rbpb = 50 rbpd = 50 rbps = 50
+ rbdb = 50 rbsb = 50 gbmin = 1E-12
+ tnom = 30 ute = -0.546000313704545 lute = -1.086399162248161E-7
+ wute = -3.970187002051872E-7 pute = 5.980103217624887E-14 kt1 = 0.051748062933343
+ lkt1 = -6.077897102454077E-8 wkt1 = -1.743576412009042E-7 pkt1 = 3.407157719480904E-14
+ kt1l = 0 kt2 = 0.047731398035249 lkt2 = -1.320766774902981E-8
+ wkt2 = -4.418592470622033E-8 pkt2 = 7.367874520430155E-15 ua1 = 2.244476856932813E-9
+ lua1 = -2.181911604389337E-16 wua1 = -5.591827841348395E-16 pua1 = 3.614327741669832E-23
+ ub1 = -2.7065105773862E-18 lub1 = 3.201682710896192E-25 wub1 = 8.059216872743307E-25
+ pub1 = -4.571496855411949E-32 uc1 = -3.723161168723502E-10 luc1 = 5.863161456792296E-17
+ wuc1 = 1.65595267031948E-16 puc1 = -1.739603382977224E-23 at = 6.318554780381558E4
+ lat = -3.803305876364924E-3 wat = -0.034452744982911 pat = 5.666834307085306E-9
+ prt = 0 njs = 1.2928 xtis = 2
+ tpb = 1.2287E-3 tpbsw = 0 tpbswg = 0
+ tcj = 7.92E-4 tcjsw = 1E-5 tcjswg = 0
+ tvoff = 0 tvfbsdoff = 0 saref = 1.75E-6
+ sbref = 1.74E-6 wlod = 0 ku0 = -2.7E-8
+ kvsat = 0.2 kvth0 = 9.8E-9 tku0 = 0
+ llodku0 = 0 wlodku0 = 1 llodvth = 0
+ wlodvth = 1 lku0 = 0 wku0 = 0
+ pku0 = 0 lkvth0 = 0 wkvth0 = 2E-7
+ pkvth0 = 0 stk2 = 0 lodk2 = 1
+ steta0 = 0 lodeta0 = 1

.model nshort_model.48 nmos
+ level = 54 lmin = 1.5E-7 lmax = 1.8E-7 wmin = 4.2E-7
+ wmax = 5.5E-7 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 4.148E-9
+ toxm = 4.148E-9 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 9.999999999999999E22 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {2.1859E-8+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {1.1932E-8-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = 0 dwb = 0 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = 0.624388294635715 lvth0 = -9.469892261755594E-9
+ wvth0 = -5.599904570804793E-9 pvth0 = -6.119141438378658E-15 k1 = -1.38213718315927
+ lk1 = 2.887518774696176E-7 wk1 = 8.613887705177163E-7 pk1 = -1.086521339580226E-13
+ k2 = 0.616568299624609 lk2 = -9.277451948795117E-8 wk2 = -2.944282428467137E-7
+ pk2 = 3.622953734046334E-14 k3 = 2 k3b = 0.54
+ w0 = 0 lpe0 = 1.0325E-7 lpeb = -7.082E-8
+ vbm = -3 dvtp0 = 0 dvtp1 = 0
+ dvt0 = 0 dvt1 = 0.53 dvt2 = -0.032
+ dvt0w = -3.58 dvt1w = 1.6706E6 dvt2w = 0.068
+ vfbsdoff = 0 u0 = 0.0935552262646 lu0 = -1.07537132179227E-8
+ wu0 = -3.725142179865745E-8 pu0 = 5.79637656634135E-15 ua = -3.081683690224791E-9
+ lua = 2.486261751703826E-16 wua = 7.7490645154577E-16 pua = -1.019390608774391E-22
+ ub = 1.100531196908236E-17 lub = -1.280647713029611E-24 wub = -4.676608354879057E-24
+ pub = 6.792941747542332E-31 uc = -3.916141613118598E-10 luc = 6.74625450104816E-17
+ wuc = 2.184857207382329E-16 puc = -3.111731619439917E-23 ud = 0
+ up = 0 lp = 1 eu = 1.67
+ vsat = 2.362930066163005E5 lvsat = -9.869301975462265E-3 wvsat = -0.034840239959817
+ pvsat = 6.068608511936989E-9 a0 = 0.888610580988553 la0 = 7.711821575642787E-8
+ wa0 = 2.300548333644653E-7 pa0 = -2.901819646126019E-14 ags = -4.54468957576923
+ lags = 7.309189643292273E-7 wags = 2.180437382949597E-6 pags = -2.750316497357303E-13
+ b0 = 0 b1 = 0 keta = -0.094248689021016
+ lketa = 3.235987291082255E-8 wketa = 4.774356241688753E-8 pketa = -1.8110875903506E-14
+ a1 = 0 a2 = 0.42385546 rdsw = 65.968
+ rdswmin = 0 rdw = 0 rdwmin = 0
+ rsw = 0 rswmin = 0 prwb = 0
+ prwg = 0.021507 wr = 1 voff = 0.130978255120153
+ lvoff = -4.269807726783563E-8 wvoff = -1.273745632531215E-7 pvoff = 1.606651791049573E-14
+ voffl = 5.8197729E-9 minv = 0 nfactor = 24.565700618111848
+ lnfactor = -2.651375197210277E-6 wnfactor = -1.086606443097673E-5 pnfactor = 1.31342459895912E-12
+ eta0 = 2.595046688830924 leta0 = -3.269878247525873E-7 weta0 = -9.764693581666778E-7
+ peta0 = 1.230396326735531E-13 etab = 0.185792236315285 letab = -2.898482124786476E-8
+ wetab = -8.6465929701188E-8 petab = 1.090646650878905E-14 dsub = -0.805056053340609
+ ldsub = 9.911624026244967E-8 wdsub = 5.376264737231109E-7 pdsub = -3.729565711843508E-14
+ cit = 0 cdsc = 0 cdscb = 0
+ cdscd = 0.019789710353989 lcdscd = -2.237363833210744E-9 wcdscd = -6.674381127419653E-9
+ pcdscd = 8.418797378882052E-16 pclm = 1.185150082225572 lpclm = -1.217273367246878E-7
+ wpclm = -3.186486268254107E-7 ppclm = 3.657015186719505E-14 pdiblc1 = -1.359264476174954
+ lpdiblc1 = 2.16479223079204E-7 wpdiblc1 = 6.457889501703641E-7 ppdiblc1 = -8.145723501868904E-14
+ pdiblc2 = -0.035883458916708 lpdiblc2 = 5.586509329763464E-9 wpdiblc2 = 1.666536836130887E-8
+ ppdiblc2 = -2.102102903622056E-15 pdiblcb = -0.05725316662666 lpdiblcb = -5.807629819099612E-9
+ wpdiblcb = -1.732500288252712E-8 ppdiblcb = 2.18530656359044E-15 drout = 3.134694447006578
+ ldrout = -3.319102071818618E-7 wdrout = -9.901363336304094E-7 pdrout = 1.248918365788053E-13
+ pscbe1 = -1.086578057994977E9 lpscbe1 = 236.88314790693437 wpscbe1 = 706.6568201046258
+ ppscbe1 = -8.913486466071707E-5 pscbe2 = 1E-12 pvag = 0
+ delta = 0.01 fprout = 0 pdits = 0
+ pditsl = 0 pditsd = 0 lambda = 0
+ vtl = 0 lc = 5E-9 xn = 3
+ alpha0 = 2.020787626948421E-5 lalpha0 = -2.54515660112766E-12 walpha0 = -7.550270798660617E-12
+ palpha0 = 9.523609574598554E-19 alpha1 = 0.85 beta0 = 27.646651014427896
+ lbeta0 = -1.740254372355877E-6 wbeta0 = -4.114326720557624E-6 pbeta0 = 5.189647152242564E-13
+ aigbacc = 1 bigbacc = 0 cigbacc = 0
+ nigbacc = 0 aigbinv = 0.35 bigbinv = 0.03
+ cigbinv = 6E-3 eigbinv = 1.1 nigbinv = 0
+ aigc = 0.43 bigc = 0.054 cigc = 0.075
+ aigsd = 0.43 bigsd = 0.054 cigsd = 0.075
+ dlcig = 0 nigc = 0 poxedge = 1
+ pigcd = 1 ntox = 1 toxref = 4.148E-9
+ agidl = 0 bgidl = 2.3E9 cgidl = 0.5
+ egidl = 0.8 noia = 2.5E42 noib = 0
+ noic = 0 em = 4.1E7 af = 1
+ ef = 0.84 kf = 0 lintnoi = -1E-7
+ tnoia = 1.5E7 tnoib = 9.9E6 ntnoi = 1
+ rnoia = 0.94 rnoib = 0.26 xpart = 0
+ cgso = {2.449068E-10/sw_func_tox_lv_ratio} cgdo = {2.449068E-10/sw_func_tox_lv_ratio} cgbo = {1E-13/sw_func_tox_lv_ratio}
+ ckappas = 0.6 cf = 1.4067E-12 clc = 1E-7
+ cle = 0.6 dlc = 9.87908E-9 dwc = 0
+ vfbcv = -1 noff = 3.4037 voffcv = -0.17287
+ acde = 0.4 moin = 6.9 cgsl = {0/sw_func_tox_lv_ratio}
+ cgdl = {0/sw_func_tox_lv_ratio} ijthsrev = 0.1 ijthsfwd = 0.1
+ xjbvs = 1 bvs = 11.7 jss = 2.75E-3
+ jsws = 6E-10 cjs = {sw_nsd_pw_cj} mjs = 0.44
+ mjsws = 9E-4 cjsws = {3.67354204E-11*sw_func_nsd_pw_cj} cjswgs = {2.38232788E-10*sw_func_nsd_pw_cj}
+ mjswgs = 0.8 pbs = 0.729 pbsws = 0.2
+ pbswgs = 0.95578 xrcrg1 = 12 xrcrg2 = 1
+ rbpb = 50 rbpd = 50 rbps = 50
+ rbdb = 50 rbsb = 50 gbmin = 1E-12
+ tnom = 30 ute = -0.748019114936554 lute = -7.709750867565507E-8
+ wute = -2.947402174798435E-7 pute = 4.383167899744458E-14 kt1 = -0.743513718991346
+ lkt1 = 6.339002255805236E-8 wkt1 = 2.282690842754882E-7 pkt1 = -2.879294921417297E-14
+ kt1l = 0 kt2 = -0.070413477856473 lkt2 = 5.239000593200037E-9
+ wkt2 = 1.562869934999126E-8 pkt2 = -1.971341621210496E-15 ua1 = 4.508682855627463E-9
+ lua1 = -5.717152282511215E-16 wua1 = -1.705509525565965E-15 pua1 = 2.151261495167885E-22
+ ub1 = -6.389620609075741E-18 lub1 = 8.952343389974977E-25 wub1 = 2.670614000338178E-24
+ pub1 = -3.368605675466564E-31 uc1 = -6.021939828686095E-10 luc1 = 9.45238250531149E-17
+ wuc1 = 2.819782927842661E-16 puc1 = -3.556761393863618E-23 at = -2.379515109001243E4
+ lat = 9.777512526121806E-3 wat = 9.584017214452739E-3 pat = -1.20888959536221E-9
+ prt = 0 njs = 1.2928 xtis = 2
+ tpb = 1.2287E-3 tpbsw = 0 tpbswg = 0
+ tcj = 7.92E-4 tcjsw = 1E-5 tcjswg = 0
+ tvoff = 0 tvfbsdoff = 0 saref = 1.1E-6
+ sbref = 1.1E-6 wlod = 0 ku0 = -2.7E-8
+ kvsat = 0.2 kvth0 = 9.8E-9 tku0 = 0
+ llodku0 = 0 wlodku0 = 1 llodvth = 0
+ wlodvth = 1 lku0 = 0 wku0 = 0
+ pku0 = 0 lkvth0 = 0 wkvth0 = 2E-7
+ pkvth0 = 0 stk2 = 0 lodk2 = 1
+ steta0 = 0 lodeta0 = 1

.ends sky130_fd_pr__nfet_01v8
