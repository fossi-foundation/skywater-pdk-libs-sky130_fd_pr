* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

******************************************************************
******************************************************************
*  *****************************************************
*  03/23/2020 Usman Suriono
*      Why     : New scalable sky130_fd_pr__pfet_01v8 5V (HV) model
*      What    : Converted from discrete phv models
*                Add process Monte Carlo
*                Replaced rsh from 1 to calculated rsh from the original model.
*                PDK netlist nrd/nrs = ratio of distance the middle of the contact to Gate.
*
*  *****************************************************
*
*  Pmos 5V (HV) Model
*  -----------------------------------------------------

.subckt  sky130_fd_pr__pfet_g5v0d10v5  d g s b  mult=1
+ 
.param  l = 1 w = 1 nf = 1 ad = 0 as = 0 pd = 0 ps = 0 nrd = {0.14/w} nrs = {0.14/w} sa = 0 sb = 0 sd = 0
+ swx_nrds = {361*nf/w+1489}

Msky130_fd_pr__pfet_g5v0d10v5  d g s b phv_model l = {l} w = {w} ad = {ad} as = {as} pd = {pd} ps = {ps} nrd = {nrd} nrs = {nrs} sa = {sa} sb = {sb} sd = {sd} nf = {nf}
* + deltox = 0.3*(sw_tox_hv_corner - sw_tox_hv_nom) + sw_tox_hv_mc + sw_mm_tox_hv * mismatch_factor*MC_MM_SWITCH*AGAUSS(0,1.0,1)/sqrt(l*w*mult)
* + mulu0  = sw_u0_sky130_fd_pr__pfet_g5v0d10v5
+ delvto = {(sw_vth0_sky130_fd_pr__pfet_g5v0d10v5+sw_vth0_sky130_fd_pr__pfet_g5v0d10v5_mc)*(0.011*8/l+0.989)*(-0.012*7/w+1.012)*(0.0030*56/(w*l)+0.9970)+sw_mm_vth0_sky130_fd_pr__pfet_g5v0d10v5*mismatch_factor*MC_MM_SWITCH*AGAUSS(0,1.0,1)/sqrt(l*w*mult)}
* + mulvsat = sw_vsat_sky130_fd_pr__pfet_g5v0d10v5




.model phv_model.1 pmos
+ level = 54 lmin = 8E-6 lmax = 2.02E-5 wmin = 2E-5
+ wmax = 1.01E-3 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 1.175E-8
+ toxm = 1.175E-8 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 1E23 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {1.2277E-8+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {4.5375E-8-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = -4.7338E-9 dwb = 0 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = -1.011028 k1 = 0.59521
+ k2 = 2.52804E-2 k3 = -2.2405 k3b = -0.172
+ w0 = 0 lpe0 = 0 lpeb = 0
+ vbm = -3 dvtp0 = 0 dvtp1 = 0
+ dvt0 = 4.657 dvt1 = 0.34864 dvt2 = -0.030206
+ dvt0w = -2.2 dvt1w = 1.0163E6 dvt2w = 0
+ vfbsdoff = 0 u0 = 2.09856E-2 ua = 2.704411E-9
+ ub = -1.7524E-19 uc = -3.9972E-11 ud = 0
+ up = 0 lp = 1 eu = 1.67
+ vsat = 2E5 a0 = 0.89674 ags = 0.134273
+ b0 = 0 b1 = 0 keta = -7.9259E-3
+ a1 = 0 a2 = 0.5 rdsw = 788.47
+ rdswmin = 0 rdw = 0 rdwmin = 0
+ rsw = 0 rswmin = 0 prwb = 0.053538
+ prwg = 0 wr = 1 voff = -9.32047E-2
+ voffl = 0 minv = 0 nfactor = 1.74009
+ eta0 = 0.08 etab = -0.07 dsub = 0.56
+ cit = 1E-5 cdsc = 0 cdscb = 0
+ cdscd = 0 pclm = 8.35312E-2 pdiblc1 = 0.39
+ pdiblc2 = 2.940788E-3 pdiblcb = -0.025 drout = 0.56
+ pscbe1 = 3.337128E8 pscbe2 = 1.500096E-8 pvag = 0
+ delta = 0.01 fprout = 0 pdits = 0
+ pditsl = 0 pditsd = 0 lambda = 0
+ vtl = 0 lc = 5E-9 xn = 3
+ alpha0 = 5.066719E-5 alpha1 = 0 beta0 = 38.266046
+ aigbacc = 0.43 bigbacc = 0.054 cigbacc = 0.075
+ nigbacc = 1 aigbinv = 0.35 bigbinv = 0.03
+ cigbinv = 6E-3 eigbinv = 1.1 nigbinv = 3
+ aigc = 0.43 bigc = 0.054 cigc = 0.075
+ aigsd = 0.43 bigsd = 0.054 cigsd = 0.075
+ dlcig = 0 nigc = 1 poxedge = 1
+ pigcd = 1 ntox = 1 toxref = 1.175E-8
+ agidl = 7.3657E-9 bgidl = 1.7047E9 cgidl = 700
+ egidl = 0.693508 noia = 3E40 noib = 8.53E24
+ noic = 8.4E7 em = 4.1E7 af = 1
+ ef = 0.88 kf = 0 lintnoi = 0
+ tnoia = 1.5 tnoib = 3.5 ntnoi = 1
+ rnoia = 0.577 rnoib = 0.37 xpart = 0
+ cgso = {1.94171E-10/sw_func_tox_hv_ratio} cgdo = {1.94171E-10/sw_func_tox_hv_ratio} cgbo = {0/sw_func_tox_hv_ratio}
+ ckappas = 0.6 cf = 1.2E-11 clc = 1E-7
+ cle = 0.6 dlc = 4.4983E-8 dwc = 0
+ vfbcv = -0.144689 noff = 4 voffcv = 0
+ acde = 0.401 moin = 15.773 cgsl = {9.82591E-12/sw_func_tox_hv_ratio}
+ cgdl = {9.82591E-12/sw_func_tox_hv_ratio} ijthsrev = 0.1 ijthsfwd = 0.1
+ xjbvs = 1 bvs = 12.69 jss = 2.1483E-5
+ jsws = 4.02E-12 cjs = {sw_psd_nw_cj} mjs = 0.33956
+ mjsws = 0.24676 cjsws = {9.960545E-11*sw_func_psd_nw_cj} cjswgs = {1.47314E-10*sw_func_psd_nw_cj}
+ mjswgs = 0.81 pbs = 0.6587 pbsws = 1
+ pbswgs = 3 xrcrg1 = 12 xrcrg2 = 1
+ rbpb = 50 rbpd = 50 rbps = 50
+ rbdb = 50 rbsb = 50 gbmin = 1E-12
+ tnom = 30 ute = -1.3864 kt1 = -0.57573
+ kt1l = 0 kt2 = -0.019032 ua1 = 7.0656E-10
+ ub1 = -3.145E-18 uc1 = -1.092E-10 at = 4.3E5
+ prt = 0 njs = 1.3632 xtis = 10
+ tpb = 1.671E-3 tpbsw = 0 tpbswg = 0
+ tcj = 9.6E-4 tcjsw = 3E-5 tcjswg = 0
+ tvoff = 0 tvfbsdoff = 0 saref = 3E-6
+ sbref = 3E-6 wlod = 0 ku0 = 7E-8
+ kvsat = 0.4 kvth0 = 3.5E-8 tku0 = 0
+ llodku0 = 0 wlodku0 = 1 llodvth = 0
+ wlodvth = 1 lku0 = 0 wku0 = 0
+ pku0 = 0 lkvth0 = 0 wkvth0 = 6.5E-7
+ pkvth0 = 0 stk2 = 0 lodk2 = 1
+ steta0 = 0 lodeta0 = 1

.model phv_model.2 pmos
+ level = 54 lmin = 4E-6 lmax = 8E-6 wmin = 2E-5
+ wmax = 1.01E-3 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 1.175E-8
+ toxm = 1.175E-8 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 1E23 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {1.2277E-8+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {4.5375E-8-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = -4.7338E-9 dwb = 0 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = -1.016266 lvth0 = 4.143178E-8
+ k1 = 0.604152 lk1 = -7.072775E-8 k2 = 2.32995E-2
+ lk2 = 1.566755E-8 k3 = -2.2405 k3b = -0.172
+ w0 = 0 lpe0 = 0 lpeb = 0
+ vbm = -3 dvtp0 = 0 dvtp1 = 0
+ dvt0 = 4.657 dvt1 = 0.34864 dvt2 = -0.030206
+ dvt0w = -2.2 dvt1w = 1.0163E6 dvt2w = 0
+ vfbsdoff = 0 u0 = 2.02516E-2 lu0 = 5.805086E-9
+ ua = 2.449766E-9 lua = 2.014057E-15 ub = 8.85171E-20
+ lub = -2.086121E-24 uc = -5.157563E-11 luc = 9.177602E-17
+ ud = 0 up = 0 lp = 1
+ eu = 1.67 vsat = 2.977215E5 lvsat = -0.772904
+ a0 = 0.916542 la0 = -1.566198E-7 ags = 0.109759
+ lags = 1.93893E-7 b0 = 0 b1 = 0
+ keta = -4.956727E-3 lketa = -2.348393E-8 a1 = 0
+ a2 = 0.5 rdsw = 788.47 rdswmin = 0
+ rdw = 0 rdwmin = 0 rsw = 0
+ rswmin = 0 prwb = 0.053538 prwg = 0
+ wr = 1 voff = -9.47765E-2 lvoff = 1.243193E-8
+ voffl = 0 minv = 0 nfactor = 1.75518
+ lnfactor = -1.193482E-7 eta0 = 0.08 etab = -0.07
+ dsub = 0.56 cit = 1E-5 cdsc = 0
+ cdscb = 0 cdscd = 0 pclm = -0.648319
+ lpclm = 5.788389E-6 pdiblc1 = 0.39 pdiblc2 = 4.554123E-3
+ lpdiblc2 = -1.276027E-8 pdiblcb = -0.025 drout = 0.56
+ pscbe1 = 5.621233E8 lpscbe1 = -1.806556E3 pscbe2 = -1.531739E-8
+ lpscbe2 = 2.397954E-13 pvag = 0 delta = 0.01
+ fprout = 0 pdits = 0 pditsl = 0
+ pditsd = 0 lambda = 0 vtl = 0
+ lc = 5E-9 xn = 3 alpha0 = 7.815322E-5
+ lalpha0 = -2.173939E-10 alpha1 = 0 beta0 = 39.140288
+ lbeta0 = -6.9146E-6 aigbacc = 0.43 bigbacc = 0.054
+ cigbacc = 0.075 nigbacc = 1 aigbinv = 0.35
+ bigbinv = 0.03 cigbinv = 6E-3 eigbinv = 1.1
+ nigbinv = 3 aigc = 0.43 bigc = 0.054
+ cigc = 0.075 aigsd = 0.43 bigsd = 0.054
+ cigsd = 0.075 dlcig = 0 nigc = 1
+ poxedge = 1 pigcd = 1 ntox = 1
+ toxref = 1.175E-8 agidl = 6.538796E-9 lagidl = 6.540191E-15
+ bgidl = 1.478354E9 lbgidl = 1.790224E3 cgidl = 932.600375
+ lcgidl = -1.839695E-3 egidl = 1.209319 legidl = -4.079675E-6
+ noia = 3E40 noib = 8.53E24 noic = 8.4E7
+ em = 4.1E7 af = 1 ef = 0.88
+ kf = 0 lintnoi = 0 tnoia = 1.5
+ tnoib = 3.5 ntnoi = 1 rnoia = 0.577
+ rnoib = 0.37 xpart = 0 cgso = {1.94171E-10/sw_func_tox_hv_ratio}
+ cgdo = {1.94171E-10/sw_func_tox_hv_ratio} cgbo = {0/sw_func_tox_hv_ratio} ckappas = 0.6
+ cf = 1.2E-11 clc = 1E-7 cle = 0.6
+ dlc = 4.4983E-8 dwc = 0 vfbcv = -0.144689
+ noff = 4 voffcv = 0 acde = 0.401
+ moin = 15.773 cgsl = {9.82591E-12/sw_func_tox_hv_ratio} cgdl = {9.82591E-12/sw_func_tox_hv_ratio}
+ ijthsrev = 0.1 ijthsfwd = 0.1 xjbvs = 1
+ bvs = 12.69 jss = 2.1483E-5 jsws = 4.02E-12
+ cjs = {sw_psd_nw_cj} mjs = 0.33956 mjsws = 0.24676
+ cjsws = {9.960545E-11*sw_func_psd_nw_cj} cjswgs = {1.47314E-10*sw_func_psd_nw_cj} mjswgs = 0.81
+ pbs = 0.6587 pbsws = 1 pbswgs = 3
+ xrcrg1 = 12 xrcrg2 = 1 rbpb = 50
+ rbpd = 50 rbps = 50 rbdb = 50
+ rbsb = 50 gbmin = 1E-12 tnom = 30
+ ute = -1.22055 lute = -1.311749E-6 kt1 = -0.585239
+ lkt1 = 7.521104E-8 kt1l = 0 kt2 = -0.019032
+ ua1 = 1.375495E-9 lua1 = -5.290776E-15 ub1 = -2.61041E-18
+ lub1 = -4.228205E-24 uc1 = -1.092E-10 at = 6.730478E5
+ lat = -1.922326 prt = 0 njs = 1.3632
+ xtis = 10 tpb = 1.671E-3 tpbsw = 0
+ tpbswg = 0 tcj = 9.6E-4 tcjsw = 3E-5
+ tcjswg = 0 tvoff = 0 tvfbsdoff = 0
+ saref = 3E-6 sbref = 3E-6 wlod = 0
+ ku0 = 7E-8 kvsat = 0.4 kvth0 = 3.5E-8
+ tku0 = 0 llodku0 = 0 wlodku0 = 1
+ llodvth = 0 wlodvth = 1 lku0 = 0
+ wku0 = 0 pku0 = 0 lkvth0 = 0
+ wkvth0 = 6.5E-7 pkvth0 = 0 stk2 = 0
+ lodk2 = 1 steta0 = 0 lodeta0 = 1

.model phv_model.3 pmos
+ level = 54 lmin = 2E-6 lmax = 4E-6 wmin = 2E-5
+ wmax = 1.01E-3 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 1.175E-8
+ toxm = 1.175E-8 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 1E23 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {1.2277E-8+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {4.5375E-8-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = -4.7338E-9 dwb = 0 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = -0.991137 lvth0 = -5.680649E-8
+ k1 = 0.602594 lk1 = -6.463595E-8 k2 = 2.68321E-2
+ lk2 = 1.857724E-9 k3 = -2.2405 k3b = -0.172
+ w0 = 0 lpe0 = 0 lpeb = 0
+ vbm = -3 dvtp0 = 0 dvtp1 = 0
+ dvt0 = 4.657 dvt1 = 0.34864 dvt2 = -0.030206
+ dvt0w = -2.2 dvt1w = 1.0163E6 dvt2w = 0
+ vfbsdoff = 0 u0 = 2.09383E-2 lu0 = 3.120588E-9
+ ua = 3.313866E-9 lua = -1.363927E-15 ub = -1.459991E-18
+ lub = 3.967386E-24 uc = -5.492301E-11 luc = 1.048618E-16
+ ud = 0 up = 0 lp = 1
+ eu = 1.67 vsat = 8.454508E4 lvsat = 6.04563E-2
+ a0 = 0.823723 la0 = 2.062331E-7 ags = 0.121307
+ lags = 1.487485E-7 b0 = 0 b1 = 0
+ keta = -5.087328E-3 lketa = -2.297338E-8 a1 = 0
+ a2 = 0.5 rdsw = 788.47 rdswmin = 0
+ rdw = 0 rdwmin = 0 rsw = 0
+ rswmin = 0 prwb = 0.053538 prwg = 0
+ wr = 1 voff = -0.064087 lvoff = -1.075408E-7
+ voffl = 0 minv = 0 nfactor = 2.156069
+ lnfactor = -1.686524E-6 eta0 = 1.90949E-2 leta0 = 2.380932E-7
+ etab = -0.122401 letab = 2.048497E-7 dsub = 0.814742
+ ldsub = -9.958489E-7 cit = 1E-5 cdsc = 0
+ cdscb = 0 cdscd = 0 pclm = 1.048766
+ lpclm = -8.459407E-7 pdiblc1 = 0.581562 lpdiblc1 = -7.488642E-7
+ pdiblc2 = -1.133342E-3 lpdiblc2 = 9.473451E-9 pdiblcb = 0.165925
+ lpdiblcb = -7.463736E-7 drout = 0.139965 ldrout = 1.642022E-6
+ pscbe1 = -1.561704E8 lpscbe1 = 1.001434E3 pscbe2 = 7.607469E-8
+ lpscbe2 = -1.174791E-13 pvag = 0 delta = 0.01
+ fprout = 0 pdits = 0 pditsl = 0
+ pditsd = 0 lambda = 0 vtl = 0
+ lc = 5E-9 xn = 3 alpha0 = 4.406319E-5
+ lalpha0 = -8.412745E-11 alpha1 = -9.54625E-11 lalpha1 = 3.731868E-16
+ beta0 = 70.183411 lbeta0 = -1.282699E-4 aigbacc = 0.43
+ bigbacc = 0.054 cigbacc = 0.075 nigbacc = 1
+ aigbinv = 0.35 bigbinv = 0.03 cigbinv = 6E-3
+ eigbinv = 1.1 nigbinv = 3 aigc = 0.43
+ bigc = 0.054 cigc = 0.075 aigsd = 0.43
+ bigsd = 0.054 cigsd = 0.075 dlcig = 0
+ nigc = 1 poxedge = 1 pigcd = 1
+ ntox = 1 toxref = 1.175E-8 agidl = 9.197164E-9
+ lagidl = -3.852034E-15 bgidl = 2.620002E9 lbgidl = -2.672764E3
+ cgidl = 455.747206 lcgidl = 2.444373E-5 egidl = -1.585323
+ legidl = 6.845277E-6 noia = 3E40 noib = 8.53E24
+ noic = 8.4E7 em = 4.1E7 af = 1
+ ef = 0.88 kf = 0 lintnoi = 0
+ tnoia = 1.5 tnoib = 3.5 ntnoi = 1
+ rnoia = 0.577 rnoib = 0.37 xpart = 0
+ cgso = {1.94171E-10/sw_func_tox_hv_ratio} cgdo = {1.94171E-10/sw_func_tox_hv_ratio} cgbo = {0/sw_func_tox_hv_ratio}
+ ckappas = 0.6 cf = 1.2E-11 clc = 1E-7
+ cle = 0.6 dlc = 4.4983E-8 dwc = 0
+ vfbcv = -0.144689 noff = 4 voffcv = 0
+ acde = 0.401 moin = 15.773 cgsl = {9.82591E-12/sw_func_tox_hv_ratio}
+ cgdl = {9.82591E-12/sw_func_tox_hv_ratio} ijthsrev = 0.1 ijthsfwd = 0.1
+ xjbvs = 1 bvs = 12.69 jss = 2.1483E-5
+ jsws = 4.02E-12 cjs = {sw_psd_nw_cj} mjs = 0.33956
+ mjsws = 0.24676 cjsws = {9.960545E-11*sw_func_psd_nw_cj} cjswgs = {1.47314E-10*sw_func_psd_nw_cj}
+ mjswgs = 0.81 pbs = 0.6587 pbsws = 1
+ pbswgs = 3 xrcrg1 = 12 xrcrg2 = 1
+ rbpb = 50 rbpd = 50 rbps = 50
+ rbdb = 50 rbsb = 50 gbmin = 1E-12
+ tnom = 30 ute = -1.705117 lute = 5.825446E-7
+ kt1 = -0.566955 lkt1 = 3.731868E-9 kt1l = 0
+ kt2 = -0.019032 ua1 = -4.841455E-10 lua1 = 1.979024E-15
+ ub1 = -3.719971E-18 lub1 = 1.093437E-25 uc1 = -1.092E-10
+ at = 2.104356E5 lat = -0.113859 prt = 0
+ njs = 1.3632 xtis = 10 tpb = 1.671E-3
+ tpbsw = 0 tpbswg = 0 tcj = 9.6E-4
+ tcjsw = 3E-5 tcjswg = 0 tvoff = 0
+ tvfbsdoff = 0 saref = 3E-6 sbref = 3E-6
+ wlod = 0 ku0 = 7E-8 kvsat = 0.4
+ kvth0 = 3.5E-8 tku0 = 0 llodku0 = 0
+ wlodku0 = 1 llodvth = 0 wlodvth = 1
+ lku0 = 0 wku0 = 0 pku0 = 0
+ lkvth0 = 0 wkvth0 = 6.5E-7 pkvth0 = 0
+ stk2 = 0 lodk2 = 1 steta0 = 0
+ lodeta0 = 1

.model phv_model.4 pmos
+ level = 54 lmin = 1E-6 lmax = 2E-6 wmin = 2E-5
+ wmax = 1.01E-3 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 1.175E-8
+ toxm = 1.175E-8 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 1E23 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {1.2277E-8+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {4.5375E-8-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = -4.7338E-9 dwb = 0 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = -1.041714 lvth0 = 3.975754E-8
+ k1 = 0.559056 lk1 = 1.848825E-8 k2 = 2.28798E-2
+ lk2 = 9.40366E-9 k3 = -2.2405 k3b = -0.172
+ w0 = 0 lpe0 = 0 lpeb = 0
+ vbm = -3 dvtp0 = 0 dvtp1 = 0
+ dvt0 = 4.657 dvt1 = 0.34864 dvt2 = -0.030206
+ dvt0w = -2.2 dvt1w = 1.0163E6 dvt2w = 0
+ vfbsdoff = 0 u0 = 2.56676E-2 lu0 = -5.908774E-9
+ ua = 3.462013E-9 lua = -1.646777E-15 ub = 4.300207E-19
+ lub = 3.588803E-25 uc = 5.323295E-13 luc = -1.01635E-18
+ ud = 0 up = 0 lp = 1
+ eu = 1.67 vsat = 1.783309E5 lvsat = -0.118604
+ a0 = 1.021774 la0 = -1.718962E-7 ags = -0.288817
+ lags = 9.317778E-7 b0 = 0 b1 = 0
+ keta = 4.43017E-2 lketa = -1.172693E-7 a1 = 0
+ a2 = 0.5 rdsw = 788.47 rdswmin = 0
+ rdw = 0 rdwmin = 0 rsw = 0
+ rswmin = 0 prwb = 0.053538 prwg = 0
+ wr = 1 voff = -0.1592 lvoff = 7.405273E-8
+ voffl = 0 minv = 0 nfactor = 1.007074
+ lnfactor = 5.071942E-7 eta0 = 0.274524 leta0 = -2.49585E-7
+ etab = -2.88449E-2 letab = 2.622727E-8 dsub = 6.49192E-2
+ ldsub = 4.357497E-7 cit = 1.454625E-5 lcit = -8.679928E-12
+ cdsc = 0 cdscb = 0 cdscd = 0
+ pclm = 6.24965E-2 lpclm = 1.037094E-6 pdiblc1 = -1.786113E-3
+ lpdiblc1 = 3.648934E-7 pdiblc2 = 5.940119E-3 lpdiblc2 = -4.031554E-9
+ pdiblcb = -0.40685 lpdiblcb = 3.471971E-7 drout = 1.535831
+ ldrout = -1.023035E-6 pscbe1 = 4.309632E8 lpscbe1 = -119.550868
+ pscbe2 = 1.454314E-8 pvag = 0 delta = 0.01
+ fprout = 0 pdits = 0 pditsl = 0
+ pditsd = 0 lambda = 0 vtl = 0
+ lc = 5E-9 xn = 3 alpha0 = -6.165893E-5
+ lalpha0 = 1.177225E-10 alpha1 = 1.90925E-10 lalpha1 = -1.735986E-16
+ beta0 = -39.873797 lbeta0 = 8.18568E-5 aigbacc = 0.43
+ bigbacc = 0.054 cigbacc = 0.075 nigbacc = 1
+ aigbinv = 0.35 bigbinv = 0.03 cigbinv = 6E-3
+ eigbinv = 1.1 nigbinv = 3 aigc = 0.43
+ bigc = 0.054 cigc = 0.075 aigsd = 0.43
+ bigsd = 0.054 cigsd = 0.075 dlcig = 0
+ nigc = 1 poxedge = 1 pigcd = 1
+ ntox = 1 toxref = 1.175E-8 agidl = 3.842289E-9
+ lagidl = 6.371761E-15 bgidl = 8.553089E8 lbgidl = 696.477408
+ cgidl = 439.517648 lcgidl = 5.543002E-5 egidl = 3.110213
+ legidl = -2.119675E-6 noia = 3E40 noib = 8.53E24
+ noic = 8.4E7 em = 4.1E7 af = 1
+ ef = 0.88 kf = 0 lintnoi = 0
+ tnoia = 1.5 tnoib = 3.5 ntnoi = 1
+ rnoia = 0.577 rnoib = 0.37 xpart = 0
+ cgso = {1.94171E-10/sw_func_tox_hv_ratio} cgdo = {1.94171E-10/sw_func_tox_hv_ratio} cgbo = {0/sw_func_tox_hv_ratio}
+ ckappas = 0.6 cf = 1.2E-11 clc = 1E-7
+ cle = 0.6 dlc = 4.4983E-8 dwc = 0
+ vfbcv = -0.144689 noff = 4 voffcv = 0
+ acde = 0.401 moin = 15.773 cgsl = {9.82591E-12/sw_func_tox_hv_ratio}
+ cgdl = {9.82591E-12/sw_func_tox_hv_ratio} ijthsrev = 0.1 ijthsfwd = 0.1
+ xjbvs = 1 bvs = 12.69 jss = 2.1483E-5
+ jsws = 4.02E-12 cjs = {sw_psd_nw_cj} mjs = 0.33956
+ mjsws = 0.24676 cjsws = {9.960545E-11*sw_func_psd_nw_cj} cjswgs = {1.47314E-10*sw_func_psd_nw_cj}
+ mjswgs = 0.81 pbs = 0.6587 pbsws = 1
+ pbswgs = 3 xrcrg1 = 12 xrcrg2 = 1
+ rbpb = 50 rbpd = 50 rbps = 50
+ rbdb = 50 rbsb = 50 gbmin = 1E-12
+ tnom = 30 ute = -1.211876 lute = -3.591754E-7
+ kt1 = -0.500261 lkt1 = -1.236022E-7 kt1l = 0
+ kt2 = -0.019032 ua1 = 6.729484E-10 lua1 = -2.30157E-16
+ ub1 = -3.532041E-18 lub1 = -2.494611E-25 uc1 = -1.092E-10
+ at = 2.608192E5 lat = -0.210054 prt = 0
+ njs = 1.3632 xtis = 10 tpb = 1.671E-3
+ tpbsw = 0 tpbswg = 0 tcj = 9.6E-4
+ tcjsw = 3E-5 tcjswg = 0 tvoff = 0
+ tvfbsdoff = 0 saref = 3E-6 sbref = 3E-6
+ wlod = 0 ku0 = 7E-8 kvsat = 0.4
+ kvth0 = 3.5E-8 tku0 = 0 llodku0 = 0
+ wlodku0 = 1 llodvth = 0 wlodvth = 1
+ lku0 = 0 wku0 = 0 pku0 = 0
+ lkvth0 = 0 wkvth0 = 6.5E-7 pkvth0 = 0
+ stk2 = 0 lodk2 = 1 steta0 = 0
+ lodeta0 = 1

.model phv_model.5 pmos
+ level = 54 lmin = 8E-7 lmax = 1E-6 wmin = 2E-5
+ wmax = 1.01E-3 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 1.175E-8
+ toxm = 1.175E-8 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 1E23 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {1.2277E-8+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {4.5375E-8-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = -4.7338E-9 dwb = 0 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = -1.086499 lvth0 = 8.047849E-8
+ k1 = 0.590242 lk1 = -9.866749E-9 k2 = 2.22322E-2
+ lk2 = 9.992502E-9 k3 = -2.2405 k3b = -0.172
+ w0 = 0 lpe0 = 0 lpeb = 0
+ vbm = -3 dvtp0 = 0 dvtp1 = 0
+ dvt0 = 4.657 dvt1 = 0.34864 dvt2 = -0.030206
+ dvt0w = -2.2 dvt1w = 1.0163E6 dvt2w = 0
+ vfbsdoff = 0 u0 = 1.91691E-2 ua = -8.205359E-10
+ lua = 2.247131E-15 ub = 4.352104E-18 lub = -3.207274E-24
+ uc = 6.082696E-12 luc = -6.063021E-18 ud = 0
+ up = 0 lp = 1 eu = 1.67
+ vsat = 8.367108E3 lvsat = 3.59353E-2 a0 = 0.794461
+ la0 = 3.478835E-8 ags = 0.788582 lags = -4.784728E-8
+ b0 = 0 b1 = 0 keta = -0.15376
+ lketa = 6.28183E-8 a1 = 0 a2 = 0.5
+ rdsw = 788.47 rdswmin = 0 rdw = 0
+ rdwmin = 0 rsw = 0 rswmin = 0
+ prwb = 0.053538 prwg = 0 wr = 1
+ voff = -9.52546E-2 lvoff = 1.591078E-8 voffl = 0
+ minv = 0 nfactor = 1.183704 lnfactor = 3.465937E-7
+ eta0 = -7.166468E-5 leta0 = 9.120294E-11 etab = 7.545356E-4
+ letab = -6.860615E-10 dsub = 1.499307 ldsub = -8.684674E-7
+ cit = -1.273125E-5 lcit = 1.612214E-11 cdsc = 0
+ cdscb = 0 cdscd = 0 pclm = 2.021902
+ lpclm = -7.444957E-7 pdiblc1 = 0.195862 lpdiblc1 = 1.851818E-7
+ pdiblc2 = -3.36185E-2 lpdiblc2 = 3.193712E-8 pdiblcb = -0.025
+ drout = 0.335842 ldrout = 6.805458E-8 pscbe1 = -5.698769E7
+ lpscbe1 = 324.118516 pscbe2 = 1.828151E-8 lpscbe2 = -3.388725E-15
+ pvag = 0 delta = 0.01 fprout = 0
+ pdits = 0 pditsl = 0 pditsd = 0
+ lambda = 0 vtl = 0 lc = 5E-9
+ xn = 3 alpha0 = 2.471576E-4 lalpha0 = -1.63069E-10
+ alpha1 = 0 beta0 = 67.196894 lbeta0 = -1.549723E-5
+ aigbacc = 0.43 bigbacc = 0.054 cigbacc = 0.075
+ nigbacc = 1 aigbinv = 0.35 bigbinv = 0.03
+ cigbinv = 6E-3 eigbinv = 1.1 nigbinv = 3
+ aigc = 0.43 bigc = 0.054 cigc = 0.075
+ aigsd = 0.43 bigsd = 0.054 cigsd = 0.075
+ dlcig = 0 nigc = 1 poxedge = 1
+ pigcd = 1 ntox = 1 toxref = 1.175E-8
+ agidl = 9.041412E-9 lagidl = 1.644458E-15 bgidl = 9.616975E8
+ lbgidl = 599.743573 cgidl = 431.2572 lcgidl = 6.294083E-5
+ egidl = 1.835557 legidl = -9.606931E-7 noia = 3E40
+ noib = 8.53E24 noic = 8.4E7 em = 4.1E7
+ af = 1 ef = 0.88 kf = 0
+ lintnoi = 0 tnoia = 1.5 tnoib = 3.5
+ ntnoi = 1 rnoia = 0.577 rnoib = 0.37
+ xpart = 0 cgso = {1.94171E-10/sw_func_tox_hv_ratio} cgdo = {1.94171E-10/sw_func_tox_hv_ratio}
+ cgbo = {0/sw_func_tox_hv_ratio} ckappas = 0.6 cf = 1.2E-11
+ clc = 1E-7 cle = 0.6 dlc = 4.4983E-8
+ dwc = 0 vfbcv = -0.144689 noff = 4
+ voffcv = 0 acde = 0.401 moin = 15.773
+ cgsl = {9.82591E-12/sw_func_tox_hv_ratio} cgdl = {9.82591E-12/sw_func_tox_hv_ratio} ijthsrev = 0.1
+ ijthsfwd = 0.1 xjbvs = 1 bvs = 12.69
+ jss = 2.1483E-5 jsws = 4.02E-12 cjs = {sw_psd_nw_cj}
+ mjs = 0.33956 mjsws = 0.24676 cjsws = {9.960545E-11*sw_func_psd_nw_cj}
+ cjswgs = {1.47314E-10*sw_func_psd_nw_cj} mjswgs = 0.81 pbs = 0.6587
+ pbsws = 1 pbswgs = 3 xrcrg1 = 12
+ xrcrg2 = 1 rbpb = 50 rbpd = 50
+ rbps = 50 rbdb = 50 rbsb = 50
+ gbmin = 1E-12 tnom = 30 ute = -2.057628
+ lute = 4.098248E-7 kt1 = -0.610312 lkt1 = -2.353832E-8
+ kt1l = 0 kt2 = -0.019032 ua1 = -5.034182E-11
+ lua1 = 4.274946E-16 ub1 = -4.570617E-18 lub1 = 6.948642E-25
+ uc1 = -1.092E-10 at = 4.6822E4 lat = -1.54773E-2
+ prt = 0 njs = 1.3632 xtis = 10
+ tpb = 1.671E-3 tpbsw = 0 tpbswg = 0
+ tcj = 9.6E-4 tcjsw = 3E-5 tcjswg = 0
+ tvoff = 0 tvfbsdoff = 0 saref = 2.81E-6
+ sbref = 2.81E-6 wlod = 0 ku0 = 7E-8
+ kvsat = 0.4 kvth0 = 3.5E-8 tku0 = 0
+ llodku0 = 0 wlodku0 = 1 llodvth = 0
+ wlodvth = 1 lku0 = 0 wku0 = 0
+ pku0 = 0 lkvth0 = 0 wkvth0 = 6.5E-7
+ pkvth0 = 0 stk2 = 0 lodk2 = 1
+ steta0 = 0 lodeta0 = 1

.model phv_model.6 pmos
+ level = 54 lmin = 6E-7 lmax = 8E-7 wmin = 2E-5
+ wmax = 1.01E-3 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 1.175E-8
+ toxm = 1.175E-8 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 1E23 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {1.2277E-8+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {4.5375E-8-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = -4.7338E-9 dwb = 0 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = -0.973029 k1 = 0.57633
+ k2 = 0.036321 k3 = -2.2405 k3b = -0.172
+ w0 = 0 lpe0 = 0 lpeb = 0
+ vbm = -3 dvtp0 = 0 dvtp1 = 0
+ dvt0 = 4.657 dvt1 = 0.34864 dvt2 = -0.030206
+ dvt0w = -2.2 dvt1w = 1.0163E6 dvt2w = 0
+ vfbsdoff = 0 u0 = 1.91724E-2 ua = 2.347784E-9
+ ub = -1.6996E-19 uc = -2.4658E-12 ud = 0
+ up = 0 lp = 1 eu = 1.67
+ vsat = 5.90337E4 a0 = 0.84351 ags = 0.72112
+ b0 = 0 b1 = 0 keta = -0.06519
+ a1 = 0 a2 = 0.5 rdsw = 788.47
+ rdswmin = 0 rdw = 0 rdwmin = 0
+ rsw = 0 rswmin = 0 prwb = 0.053538
+ prwg = 0 wr = 1 voff = -7.28213E-2
+ voffl = 0 minv = 0 nfactor = 1.67238
+ eta0 = 5.6926E-5 etab = -2.1277E-4 dsub = 0.27482
+ cit = 1E-5 cdsc = 0 cdscb = 0
+ cdscd = 0 pclm = 0.972208 pdiblc1 = 0.456957
+ pdiblc2 = 1.14109E-2 pdiblcb = -0.025 drout = 0.431795
+ pscbe1 = 4E8 pscbe2 = 1.350362E-8 pvag = 0
+ delta = 0.01 fprout = 0 pdits = 0
+ pditsl = 0 pditsd = 0 lambda = 0
+ vtl = 0 lc = 5E-9 xn = 3
+ alpha0 = 1.724017E-5 alpha1 = 0 beta0 = 45.34673
+ aigbacc = 0.43 bigbacc = 0.054 cigbacc = 0.075
+ nigbacc = 1 aigbinv = 0.35 bigbinv = 0.03
+ cigbinv = 6E-3 eigbinv = 1.1 nigbinv = 3
+ aigc = 0.43 bigc = 0.054 cigc = 0.075
+ aigsd = 0.43 bigsd = 0.054 cigsd = 0.075
+ dlcig = 0 nigc = 1 poxedge = 1
+ pigcd = 1 ntox = 1 toxref = 1.175E-8
+ agidl = 1.136E-8 bgidl = 1.8073E9 cgidl = 520
+ egidl = 0.481037 noia = 3E40 noib = 8.53E24
+ noic = 8.4E7 em = 4.1E7 af = 1
+ ef = 0.88 kf = 0 lintnoi = 0
+ tnoia = 1.5 tnoib = 3.5 ntnoi = 1
+ rnoia = 0.577 rnoib = 0.37 xpart = 0
+ cgso = {1.94171E-10/sw_func_tox_hv_ratio} cgdo = {1.94171E-10/sw_func_tox_hv_ratio} cgbo = {0/sw_func_tox_hv_ratio}
+ ckappas = 0.6 cf = 1.2E-11 clc = 1E-7
+ cle = 0.6 dlc = 4.4983E-8 dwc = 0
+ vfbcv = -0.144689 noff = 4 voffcv = 0
+ acde = 0.401 moin = 15.773 cgsl = {9.82591E-12/sw_func_tox_hv_ratio}
+ cgdl = {9.82591E-12/sw_func_tox_hv_ratio} ijthsrev = 0.1 ijthsfwd = 0.1
+ xjbvs = 1 bvs = 12.69 jss = 2.1483E-5
+ jsws = 4.02E-12 cjs = {sw_psd_nw_cj} mjs = 0.33956
+ mjsws = 0.24676 cjsws = {9.960545E-11*sw_func_psd_nw_cj} cjswgs = {1.47314E-10*sw_func_psd_nw_cj}
+ mjswgs = 0.81 pbs = 0.6587 pbsws = 1
+ pbswgs = 3 xrcrg1 = 12 xrcrg2 = 1
+ rbpb = 50 rbpd = 50 rbps = 50
+ rbdb = 50 rbsb = 50 gbmin = 1E-12
+ tnom = 30 ute = -1.4798 kt1 = -0.6435
+ kt1l = 0 kt2 = -0.019032 ua1 = 5.524E-10
+ ub1 = -3.5909E-18 uc1 = -1.092E-10 at = 2.5E4
+ prt = 0 njs = 1.3632 xtis = 10
+ tpb = 1.671E-3 tpbsw = 0 tpbswg = 0
+ tcj = 9.6E-4 tcjsw = 3E-5 tcjswg = 0
+ tvoff = 0 tvfbsdoff = 0 saref = 2.41E-6
+ sbref = 2.41E-6 wlod = 0 ku0 = 7E-8
+ kvsat = 0.4 kvth0 = 3.5E-8 tku0 = 0
+ llodku0 = 0 wlodku0 = 1 llodvth = 0
+ wlodvth = 1 lku0 = 0 wku0 = 0
+ pku0 = 0 lkvth0 = 0 wkvth0 = 6.5E-7
+ pkvth0 = 0 stk2 = 0 lodk2 = 1
+ steta0 = 0 lodeta0 = 1

.model phv_model.7 pmos
+ level = 54 lmin = 5E-7 lmax = 6E-7 wmin = 2E-5
+ wmax = 1.01E-3 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 1.175E-8
+ toxm = 1.175E-8 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 1E23 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {1.2277E-8+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {4.5375E-8-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = -4.7338E-9 dwb = 0 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = -0.783264 lvth0 = -9.663789E-8
+ k1 = 0.487482 lk1 = 4.524593E-8 k2 = 2.82588E-2
+ lk2 = 4.105688E-9 k3 = -2.2405 k3b = -0.172
+ w0 = 0 lpe0 = 0 lpeb = 0
+ vbm = -3 dvtp0 = 0 dvtp1 = 0
+ dvt0 = 4.657 dvt1 = 0.34864 dvt2 = -0.030206
+ dvt0w = -2.2 dvt1w = 1.0163E6 dvt2w = 0
+ vfbsdoff = 0 u0 = 1.31838E-2 lu0 = 3.049672E-9
+ ua = 3.115935E-9 lua = -3.911812E-16 ub = -3.240604E-18
+ lub = 1.563725E-24 uc = 9.057452E-12 luc = -5.868216E-18
+ ud = 0 up = 0 lp = 1
+ eu = 1.67 vsat = 4.293708E4 lvsat = 8.197204E-3
+ a0 = 0.368248 la0 = 2.420272E-7 ags = -1.443321
+ lags = 1.102242E-6 b0 = 0 b1 = 0
+ keta = 1.94429E-2 lketa = -4.30993E-8 a1 = 0
+ a2 = 0.5 rdsw = 788.47 rdswmin = 0
+ rdw = 0 rdwmin = 0 rsw = 0
+ rswmin = 0 prwb = 0.053538 prwg = 0
+ wr = 1 voff = 4.46966E-2 lvoff = -5.984601E-8
+ voffl = 0 minv = 0 nfactor = 1.690346
+ lnfactor = -9.149224E-9 eta0 = -0.327335 leta0 = 1.667244E-7
+ etab = 1.46738E-2 letab = -7.580997E-9 dsub = 0.254971
+ ldsub = 1.010791E-8 cit = 3.04625E-5 lcit = -1.042053E-11
+ cdsc = 0 cdscb = 0 cdscd = 0
+ pclm = -0.519068 lpclm = 7.594321E-7 pdiblc1 = 1.123736
+ lpdiblc1 = -3.39557E-7 pdiblc2 = 3.84625E-2 lpdiblc2 = -1.377603E-8
+ pdiblcb = -0.025 drout = -1.482714 ldrout = 9.749638E-7
+ pscbe1 = 5.52896E8 lpscbe1 = -77.86227 pscbe2 = 9.480217E-9
+ lpscbe2 = 2.048916E-15 pvag = 0 delta = 0.01
+ fprout = 0 pdits = 0 pditsl = 0
+ pditsd = 0 lambda = 0 vtl = 0
+ lc = 5E-9 xn = 3 alpha0 = -3.097308E-4
+ lalpha0 = 1.6651E-10 alpha1 = 0 beta0 = 7.131861
+ lbeta0 = 1.946092E-5 aigbacc = 0.43 bigbacc = 0.054
+ cigbacc = 0.075 nigbacc = 1 aigbinv = 0.35
+ bigbinv = 0.03 cigbinv = 6E-3 eigbinv = 1.1
+ nigbinv = 3 aigc = 0.43 bigc = 0.054
+ cigc = 0.075 aigsd = 0.43 bigsd = 0.054
+ cigsd = 0.075 dlcig = 0 nigc = 1
+ poxedge = 1 pigcd = 1 ntox = 1
+ toxref = 1.175E-8 agidl = 1.01416E-9 lagidl = 5.268619E-15
+ bgidl = 2.596334E9 lbgidl = -401.815565 cgidl = -936.93
+ lcgidl = 7.419416E-4 egidl = -0.272932 legidl = 3.839585E-7
+ noia = 3E40 noib = 8.53E24 noic = 8.4E7
+ em = 4.1E7 af = 1 ef = 0.88
+ kf = 0 lintnoi = 0 tnoia = 1.5
+ tnoib = 3.5 ntnoi = 1 rnoia = 0.577
+ rnoib = 0.37 xpart = 0 cgso = {1.94171E-10/sw_func_tox_hv_ratio}
+ cgdo = {1.94171E-10/sw_func_tox_hv_ratio} cgbo = {0/sw_func_tox_hv_ratio} ckappas = 0.6
+ cf = 1.2E-11 clc = 1E-7 cle = 0.6
+ dlc = 4.4983E-8 dwc = 0 vfbcv = -0.144689
+ noff = 4 voffcv = 0 acde = 0.401
+ moin = 15.773 cgsl = {9.82591E-12/sw_func_tox_hv_ratio} cgdl = {9.82591E-12/sw_func_tox_hv_ratio}
+ ijthsrev = 0.1 ijthsfwd = 0.1 xjbvs = 1
+ bvs = 12.69 jss = 2.1483E-5 jsws = 4.02E-12
+ cjs = {sw_psd_nw_cj} mjs = 0.33956 mjsws = 0.24676
+ cjsws = {9.960545E-11*sw_func_psd_nw_cj} cjswgs = {1.47314E-10*sw_func_psd_nw_cj} mjswgs = 0.81
+ pbs = 0.6587 pbsws = 1 pbswgs = 3
+ xrcrg1 = 12 xrcrg2 = 1 rbpb = 50
+ rbpd = 50 rbps = 50 rbdb = 50
+ rbsb = 50 gbmin = 1E-12 tnom = 30
+ ute = -1.919334 lute = 2.238329E-7 kt1 = -0.766357
+ lkt1 = 6.256485E-8 kt1l = 0 kt2 = -0.019032
+ ua1 = 5.524E-10 ub1 = -9.446858E-18 lub1 = 2.982147E-24
+ uc1 = -3.862786E-10 luc1 = 1.411023E-16 at = 5.36475E4
+ lat = -1.45887E-2 prt = 0 njs = 1.3632
+ xtis = 10 tpb = 1.671E-3 tpbsw = 0
+ tpbswg = 0 tcj = 9.6E-4 tcjsw = 3E-5
+ tcjswg = 0 tvoff = 0 tvfbsdoff = 0
+ saref = 2.41E-6 sbref = 2.41E-6 wlod = 0
+ ku0 = 7E-8 kvsat = 0.4 kvth0 = 3.5E-8
+ tku0 = 0 llodku0 = 0 wlodku0 = 1
+ llodvth = 0 wlodvth = 1 lku0 = 0
+ wku0 = 0 pku0 = 0 lkvth0 = 0
+ wkvth0 = 6.5E-7 pkvth0 = 0 stk2 = 0
+ lodk2 = 1 steta0 = 0 lodeta0 = 1

.model phv_model.8 pmos
+ level = 54 lmin = 8E-6 lmax = 2.02E-5 wmin = 1.5E-5
+ wmax = 2E-5 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 1.175E-8
+ toxm = 1.175E-8 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 1E23 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {1.2277E-8+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {4.5375E-8-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = -4.7338E-9 dwb = 0 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = -1.011028 k1 = 0.59521
+ k2 = 2.52804E-2 k3 = -2.2405 k3b = -0.172
+ w0 = 0 lpe0 = 0 lpeb = 0
+ vbm = -3 dvtp0 = 0 dvtp1 = 0
+ dvt0 = 4.657 dvt1 = 0.34864 dvt2 = -0.030206
+ dvt0w = -2.2 dvt1w = 1.0163E6 dvt2w = 0
+ vfbsdoff = 0 u0 = 2.09856E-2 ua = 2.704411E-9
+ ub = -1.7524E-19 uc = -3.9972E-11 ud = 0
+ up = 0 lp = 1 eu = 1.67
+ vsat = 2E5 a0 = 0.89674 ags = 0.134273
+ b0 = 0 b1 = 0 keta = -7.9259E-3
+ a1 = 0 a2 = 0.5 rdsw = 788.47
+ rdswmin = 0 rdw = 0 rdwmin = 0
+ rsw = 0 rswmin = 0 prwb = 0.053538
+ prwg = 0 wr = 1 voff = -9.32047E-2
+ voffl = 0 minv = 0 nfactor = 1.74009
+ eta0 = 0.08 etab = -0.07 dsub = 0.56
+ cit = 1E-5 cdsc = 0 cdscb = 0
+ cdscd = 0 pclm = 8.35312E-2 pdiblc1 = 0.39
+ pdiblc2 = 2.940788E-3 pdiblcb = -0.025 drout = 0.56
+ pscbe1 = 3.337128E8 pscbe2 = 1.500096E-8 pvag = 0
+ delta = 0.01 fprout = 0 pdits = 0
+ pditsl = 0 pditsd = 0 lambda = 0
+ vtl = 0 lc = 5E-9 xn = 3
+ alpha0 = 5.066719E-5 alpha1 = 0 beta0 = 38.266046
+ aigbacc = 0.43 bigbacc = 0.054 cigbacc = 0.075
+ nigbacc = 1 aigbinv = 0.35 bigbinv = 0.03
+ cigbinv = 6E-3 eigbinv = 1.1 nigbinv = 3
+ aigc = 0.43 bigc = 0.054 cigc = 0.075
+ aigsd = 0.43 bigsd = 0.054 cigsd = 0.075
+ dlcig = 0 nigc = 1 poxedge = 1
+ pigcd = 1 ntox = 1 toxref = 1.175E-8
+ agidl = 7.3657E-9 bgidl = 1.7047E9 cgidl = 700
+ egidl = 0.693508 noia = 3E40 noib = 8.53E24
+ noic = 8.4E7 em = 4.1E7 af = 1
+ ef = 0.88 kf = 0 lintnoi = 0
+ tnoia = 1.5 tnoib = 3.5 ntnoi = 1
+ rnoia = 0.577 rnoib = 0.37 xpart = 0
+ cgso = {1.94171E-10/sw_func_tox_hv_ratio} cgdo = {1.94171E-10/sw_func_tox_hv_ratio} cgbo = {0/sw_func_tox_hv_ratio}
+ ckappas = 0.6 cf = 1.2E-11 clc = 1E-7
+ cle = 0.6 dlc = 4.4983E-8 dwc = 0
+ vfbcv = -0.144689 noff = 4 voffcv = 0
+ acde = 0.401 moin = 15.773 cgsl = {9.82591E-12/sw_func_tox_hv_ratio}
+ cgdl = {9.82591E-12/sw_func_tox_hv_ratio} ijthsrev = 0.1 ijthsfwd = 0.1
+ xjbvs = 1 bvs = 12.69 jss = 2.1483E-5
+ jsws = 4.02E-12 cjs = {sw_psd_nw_cj} mjs = 0.33956
+ mjsws = 0.24676 cjsws = {9.960545E-11*sw_func_psd_nw_cj} cjswgs = {1.47314E-10*sw_func_psd_nw_cj}
+ mjswgs = 0.81 pbs = 0.6587 pbsws = 1
+ pbswgs = 3 xrcrg1 = 12 xrcrg2 = 1
+ rbpb = 50 rbpd = 50 rbps = 50
+ rbdb = 50 rbsb = 50 gbmin = 1E-12
+ tnom = 30 ute = -1.3864 kt1 = -0.57573
+ kt1l = 0 kt2 = -0.019032 ua1 = 7.0656E-10
+ ub1 = -3.145E-18 uc1 = -1.092E-10 at = 4.3E5
+ prt = 0 njs = 1.3632 xtis = 10
+ tpb = 1.671E-3 tpbsw = 0 tpbswg = 0
+ tcj = 9.6E-4 tcjsw = 3E-5 tcjswg = 0
+ tvoff = 0 tvfbsdoff = 0 saref = 3E-6
+ sbref = 3E-6 wlod = 0 ku0 = 7E-8
+ kvsat = 0.4 kvth0 = 3.5E-8 tku0 = 0
+ llodku0 = 0 wlodku0 = 1 llodvth = 0
+ wlodvth = 1 lku0 = 0 wku0 = 0
+ pku0 = 0 lkvth0 = 0 wkvth0 = 6.5E-7
+ pkvth0 = 0 stk2 = 0 lodk2 = 1
+ steta0 = 0 lodeta0 = 1

.model phv_model.9 pmos
+ level = 54 lmin = 4E-6 lmax = 8E-6 wmin = 1.5E-5
+ wmax = 2E-5 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 1.175E-8
+ toxm = 1.175E-8 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 1E23 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {1.2277E-8+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {4.5375E-8-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = -4.7338E-9 dwb = 0 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = -1.016266 lvth0 = 4.143178E-8
+ k1 = 0.604152 lk1 = -7.072775E-8 k2 = 2.32995E-2
+ lk2 = 1.566755E-8 k3 = -2.2405 k3b = -0.172
+ w0 = 0 lpe0 = 0 lpeb = 0
+ vbm = -3 dvtp0 = 0 dvtp1 = 0
+ dvt0 = 4.657 dvt1 = 0.34864 dvt2 = -0.030206
+ dvt0w = -2.2 dvt1w = 1.0163E6 dvt2w = 0
+ vfbsdoff = 0 u0 = 2.02516E-2 lu0 = 5.805086E-9
+ ua = 2.449766E-9 lua = 2.014057E-15 ub = 8.85171E-20
+ lub = -2.086121E-24 uc = -5.157563E-11 luc = 9.177602E-17
+ ud = 0 up = 0 lp = 1
+ eu = 1.67 vsat = 2.977215E5 lvsat = -0.772904
+ a0 = 0.916542 la0 = -1.566198E-7 ags = 0.109759
+ lags = 1.93893E-7 b0 = 0 b1 = 0
+ keta = -4.956727E-3 lketa = -2.348393E-8 a1 = 0
+ a2 = 0.5 rdsw = 788.47 rdswmin = 0
+ rdw = 0 rdwmin = 0 rsw = 0
+ rswmin = 0 prwb = 0.053538 prwg = 0
+ wr = 1 voff = -9.47765E-2 lvoff = 1.243193E-8
+ voffl = 0 minv = 0 nfactor = 1.75518
+ lnfactor = -1.193482E-7 eta0 = 0.08 etab = -0.07
+ dsub = 0.56 cit = 1E-5 cdsc = 0
+ cdscb = 0 cdscd = 0 pclm = -0.648319
+ lpclm = 5.788389E-6 pdiblc1 = 0.39 pdiblc2 = 4.554123E-3
+ lpdiblc2 = -1.276027E-8 pdiblcb = -0.025 drout = 0.56
+ pscbe1 = 5.621233E8 lpscbe1 = -1.806556E3 pscbe2 = -1.531739E-8
+ lpscbe2 = 2.397954E-13 pvag = 0 delta = 0.01
+ fprout = 0 pdits = 0 pditsl = 0
+ pditsd = 0 lambda = 0 vtl = 0
+ lc = 5E-9 xn = 3 alpha0 = 7.815322E-5
+ lalpha0 = -2.173939E-10 alpha1 = 0 beta0 = 39.140288
+ lbeta0 = -6.9146E-6 aigbacc = 0.43 bigbacc = 0.054
+ cigbacc = 0.075 nigbacc = 1 aigbinv = 0.35
+ bigbinv = 0.03 cigbinv = 6E-3 eigbinv = 1.1
+ nigbinv = 3 aigc = 0.43 bigc = 0.054
+ cigc = 0.075 aigsd = 0.43 bigsd = 0.054
+ cigsd = 0.075 dlcig = 0 nigc = 1
+ poxedge = 1 pigcd = 1 ntox = 1
+ toxref = 1.175E-8 agidl = 6.538796E-9 lagidl = 6.540191E-15
+ bgidl = 1.478354E9 lbgidl = 1.790224E3 cgidl = 932.600375
+ lcgidl = -1.839695E-3 egidl = 1.209319 legidl = -4.079675E-6
+ noia = 3E40 noib = 8.53E24 noic = 8.4E7
+ em = 4.1E7 af = 1 ef = 0.88
+ kf = 0 lintnoi = 0 tnoia = 1.5
+ tnoib = 3.5 ntnoi = 1 rnoia = 0.577
+ rnoib = 0.37 xpart = 0 cgso = {1.94171E-10/sw_func_tox_hv_ratio}
+ cgdo = {1.94171E-10/sw_func_tox_hv_ratio} cgbo = {0/sw_func_tox_hv_ratio} ckappas = 0.6
+ cf = 1.2E-11 clc = 1E-7 cle = 0.6
+ dlc = 4.4983E-8 dwc = 0 vfbcv = -0.144689
+ noff = 4 voffcv = 0 acde = 0.401
+ moin = 15.773 cgsl = {9.82591E-12/sw_func_tox_hv_ratio} cgdl = {9.82591E-12/sw_func_tox_hv_ratio}
+ ijthsrev = 0.1 ijthsfwd = 0.1 xjbvs = 1
+ bvs = 12.69 jss = 2.1483E-5 jsws = 4.02E-12
+ cjs = {sw_psd_nw_cj} mjs = 0.33956 mjsws = 0.24676
+ cjsws = {9.960545E-11*sw_func_psd_nw_cj} cjswgs = {1.47314E-10*sw_func_psd_nw_cj} mjswgs = 0.81
+ pbs = 0.6587 pbsws = 1 pbswgs = 3
+ xrcrg1 = 12 xrcrg2 = 1 rbpb = 50
+ rbpd = 50 rbps = 50 rbdb = 50
+ rbsb = 50 gbmin = 1E-12 tnom = 30
+ ute = -1.22055 lute = -1.311749E-6 kt1 = -0.585239
+ lkt1 = 7.521104E-8 kt1l = 0 kt2 = -0.019032
+ ua1 = 1.375495E-9 lua1 = -5.290776E-15 ub1 = -2.61041E-18
+ lub1 = -4.228205E-24 uc1 = -1.092E-10 at = 6.730478E5
+ lat = -1.922326 prt = 0 njs = 1.3632
+ xtis = 10 tpb = 1.671E-3 tpbsw = 0
+ tpbswg = 0 tcj = 9.6E-4 tcjsw = 3E-5
+ tcjswg = 0 tvoff = 0 tvfbsdoff = 0
+ saref = 3E-6 sbref = 3E-6 wlod = 0
+ ku0 = 7E-8 kvsat = 0.4 kvth0 = 3.5E-8
+ tku0 = 0 llodku0 = 0 wlodku0 = 1
+ llodvth = 0 wlodvth = 1 lku0 = 0
+ wku0 = 0 pku0 = 0 lkvth0 = 0
+ wkvth0 = 6.5E-7 pkvth0 = 0 stk2 = 0
+ lodk2 = 1 steta0 = 0 lodeta0 = 1

.model phv_model.10 pmos
+ level = 54 lmin = 2E-6 lmax = 4E-6 wmin = 1.5E-5
+ wmax = 2E-5 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 1.175E-8
+ toxm = 1.175E-8 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 1E23 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {1.2277E-8+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {4.5375E-8-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = -4.7338E-9 dwb = 0 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = -0.991137 lvth0 = -5.680649E-8
+ k1 = 0.602594 lk1 = -6.463595E-8 k2 = 2.68321E-2
+ lk2 = 1.857724E-9 k3 = -2.2405 k3b = -0.172
+ w0 = 0 lpe0 = 0 lpeb = 0
+ vbm = -3 dvtp0 = 0 dvtp1 = 0
+ dvt0 = 4.657 dvt1 = 0.34864 dvt2 = -0.030206
+ dvt0w = -2.2 dvt1w = 1.0163E6 dvt2w = 0
+ vfbsdoff = 0 u0 = 2.09383E-2 lu0 = 3.120588E-9
+ ua = 3.313866E-9 lua = -1.363927E-15 ub = -1.459991E-18
+ lub = 3.967386E-24 uc = -5.492301E-11 luc = 1.048618E-16
+ ud = 0 up = 0 lp = 1
+ eu = 1.67 vsat = 8.454508E4 lvsat = 6.04563E-2
+ a0 = 0.823723 la0 = 2.062331E-7 ags = 0.121307
+ lags = 1.487485E-7 b0 = 0 b1 = 0
+ keta = -5.087328E-3 lketa = -2.297338E-8 a1 = 0
+ a2 = 0.5 rdsw = 788.47 rdswmin = 0
+ rdw = 0 rdwmin = 0 rsw = 0
+ rswmin = 0 prwb = 0.053538 prwg = 0
+ wr = 1 voff = -0.064087 lvoff = -1.075408E-7
+ voffl = 0 minv = 0 nfactor = 2.156069
+ lnfactor = -1.686524E-6 eta0 = 1.90949E-2 leta0 = 2.380932E-7
+ etab = -0.122401 letab = 2.048497E-7 dsub = 0.814742
+ ldsub = -9.958489E-7 cit = 1E-5 cdsc = 0
+ cdscb = 0 cdscd = 0 pclm = 1.048766
+ lpclm = -8.459407E-7 pdiblc1 = 0.581562 lpdiblc1 = -7.488642E-7
+ pdiblc2 = -1.133342E-3 lpdiblc2 = 9.473451E-9 pdiblcb = 0.165925
+ lpdiblcb = -7.463736E-7 drout = 0.139965 ldrout = 1.642022E-6
+ pscbe1 = -1.561704E8 lpscbe1 = 1.001434E3 pscbe2 = 7.607469E-8
+ lpscbe2 = -1.174791E-13 pvag = 0 delta = 0.01
+ fprout = 0 pdits = 0 pditsl = 0
+ pditsd = 0 lambda = 0 vtl = 0
+ lc = 5E-9 xn = 3 alpha0 = 4.406319E-5
+ lalpha0 = -8.412745E-11 alpha1 = -9.54625E-11 lalpha1 = 3.731868E-16
+ beta0 = 70.183411 lbeta0 = -1.282699E-4 aigbacc = 0.43
+ bigbacc = 0.054 cigbacc = 0.075 nigbacc = 1
+ aigbinv = 0.35 bigbinv = 0.03 cigbinv = 6E-3
+ eigbinv = 1.1 nigbinv = 3 aigc = 0.43
+ bigc = 0.054 cigc = 0.075 aigsd = 0.43
+ bigsd = 0.054 cigsd = 0.075 dlcig = 0
+ nigc = 1 poxedge = 1 pigcd = 1
+ ntox = 1 toxref = 1.175E-8 agidl = 9.197164E-9
+ lagidl = -3.852034E-15 bgidl = 2.620002E9 lbgidl = -2.672764E3
+ cgidl = 455.747206 lcgidl = 2.444373E-5 egidl = -1.585323
+ legidl = 6.845277E-6 noia = 3E40 noib = 8.53E24
+ noic = 8.4E7 em = 4.1E7 af = 1
+ ef = 0.88 kf = 0 lintnoi = 0
+ tnoia = 1.5 tnoib = 3.5 ntnoi = 1
+ rnoia = 0.577 rnoib = 0.37 xpart = 0
+ cgso = {1.94171E-10/sw_func_tox_hv_ratio} cgdo = {1.94171E-10/sw_func_tox_hv_ratio} cgbo = {0/sw_func_tox_hv_ratio}
+ ckappas = 0.6 cf = 1.2E-11 clc = 1E-7
+ cle = 0.6 dlc = 4.4983E-8 dwc = 0
+ vfbcv = -0.144689 noff = 4 voffcv = 0
+ acde = 0.401 moin = 15.773 cgsl = {9.82591E-12/sw_func_tox_hv_ratio}
+ cgdl = {9.82591E-12/sw_func_tox_hv_ratio} ijthsrev = 0.1 ijthsfwd = 0.1
+ xjbvs = 1 bvs = 12.69 jss = 2.1483E-5
+ jsws = 4.02E-12 cjs = {sw_psd_nw_cj} mjs = 0.33956
+ mjsws = 0.24676 cjsws = {9.960545E-11*sw_func_psd_nw_cj} cjswgs = {1.47314E-10*sw_func_psd_nw_cj}
+ mjswgs = 0.81 pbs = 0.6587 pbsws = 1
+ pbswgs = 3 xrcrg1 = 12 xrcrg2 = 1
+ rbpb = 50 rbpd = 50 rbps = 50
+ rbdb = 50 rbsb = 50 gbmin = 1E-12
+ tnom = 30 ute = -1.705117 lute = 5.825446E-7
+ kt1 = -0.566955 lkt1 = 3.731868E-9 kt1l = 0
+ kt2 = -0.019032 ua1 = -4.841455E-10 lua1 = 1.979024E-15
+ ub1 = -3.719971E-18 lub1 = 1.093437E-25 uc1 = -1.092E-10
+ at = 2.104356E5 lat = -0.113859 prt = 0
+ njs = 1.3632 xtis = 10 tpb = 1.671E-3
+ tpbsw = 0 tpbswg = 0 tcj = 9.6E-4
+ tcjsw = 3E-5 tcjswg = 0 tvoff = 0
+ tvfbsdoff = 0 saref = 3E-6 sbref = 3E-6
+ wlod = 0 ku0 = 7E-8 kvsat = 0.4
+ kvth0 = 3.5E-8 tku0 = 0 llodku0 = 0
+ wlodku0 = 1 llodvth = 0 wlodvth = 1
+ lku0 = 0 wku0 = 0 pku0 = 0
+ lkvth0 = 0 wkvth0 = 6.5E-7 pkvth0 = 0
+ stk2 = 0 lodk2 = 1 steta0 = 0
+ lodeta0 = 1

.model phv_model.11 pmos
+ level = 54 lmin = 1E-6 lmax = 2E-6 wmin = 1.5E-5
+ wmax = 2E-5 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 1.175E-8
+ toxm = 1.175E-8 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 1E23 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {1.2277E-8+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {4.5375E-8-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = -4.7338E-9 dwb = 0 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = -1.031624 lvth0 = 2.049365E-8
+ wvth0 = -2.015477E-7 pvth0 = 3.848049E-13 k1 = 0.559056
+ lk1 = 1.848825E-8 k2 = 2.32556E-2 lk2 = 8.686139E-9
+ wk2 = -7.507038E-9 pk2 = 1.433281E-14 k3 = -2.2405
+ k3b = -0.172 w0 = 0 lpe0 = 0
+ lpeb = 0 vbm = -3 dvtp0 = 0
+ dvtp1 = 0 dvt0 = 4.657 dvt1 = 0.34864
+ dvt2 = -0.030206 dvt0w = -2.2 dvt1w = 1.0163E6
+ dvt2w = 0 vfbsdoff = 0 u0 = 2.51605E-2
+ lu0 = -4.94064E-9 wu0 = 1.012906E-8 pu0 = -1.933891E-14
+ ua = 3.459918E-9 lua = -1.642778E-15 wua = 4.184412E-17
+ pua = -7.989089E-23 ub = 3.46307E-19 lub = 5.187108E-25
+ wub = 1.67222E-24 pub = -3.192686E-30 uc = 5.323295E-13
+ luc = -1.01635E-18 ud = 0 up = 0
+ lp = 1 eu = 1.67 vsat = 1.783309E5
+ lvsat = -0.118604 a0 = 1.021093 la0 = -1.705964E-7
+ wa0 = 1.359971E-8 pa0 = -2.596524E-14 ags = -0.284887
+ lags = 9.24275E-7 wags = -7.849751E-8 pags = 1.498714E-13
+ b0 = 0 b1 = 0 keta = 4.43017E-2
+ lketa = -1.172693E-7 a1 = 0 a2 = 0.5
+ rdsw = 788.47 rdswmin = 0 rdw = 0
+ rdwmin = 0 rsw = 0 rswmin = 0
+ prwb = 0.053538 prwg = 0 wr = 1
+ voff = -0.1592 lvoff = 7.405273E-8 voffl = 0
+ minv = 0 nfactor = 1.087983 lnfactor = 3.527191E-7
+ wnfactor = -1.616189E-6 pnfactor = 3.085709E-12 eta0 = 0.274561
+ leta0 = -2.496551E-7 weta0 = -7.331874E-10 peta0 = 1.399838E-15
+ etab = -2.88449E-2 letab = 2.622727E-8 dsub = 6.49192E-2
+ ldsub = 4.357497E-7 cit = 1.454625E-5 lcit = -8.679928E-12
+ cdsc = 0 cdscb = 0 cdscd = 0
+ pclm = 6.24965E-2 lpclm = 1.037094E-6 pdiblc1 = -1.786113E-3
+ lpdiblc1 = 3.648934E-7 pdiblc2 = 5.940119E-3 lpdiblc2 = -4.031554E-9
+ pdiblcb = -0.40685 lpdiblcb = 3.471971E-7 drout = 1.535831
+ ldrout = -1.023035E-6 pscbe1 = 4.309632E8 lpscbe1 = -119.550868
+ pscbe2 = 1.454314E-8 pvag = 0 delta = 0.01
+ fprout = 0 pdits = 0 pditsl = 0
+ pditsd = 0 lambda = 0 vtl = 0
+ lc = 5E-9 xn = 3 alpha0 = -6.165893E-5
+ lalpha0 = 1.177225E-10 alpha1 = 1.90925E-10 lalpha1 = -1.735986E-16
+ beta0 = -39.873797 lbeta0 = 8.18568E-5 aigbacc = 0.43
+ bigbacc = 0.054 cigbacc = 0.075 nigbacc = 1
+ aigbinv = 0.35 bigbinv = 0.03 cigbinv = 6E-3
+ eigbinv = 1.1 nigbinv = 3 aigc = 0.43
+ bigc = 0.054 cigc = 0.075 aigsd = 0.43
+ bigsd = 0.054 cigsd = 0.075 dlcig = 0
+ nigc = 1 poxedge = 1 pigcd = 1
+ ntox = 1 toxref = 1.175E-8 agidl = -2.975727E-9
+ lagidl = 1.938906E-14 wagidl = 1.361929E-13 pagidl = -2.600263E-19
+ bgidl = 1.039403E9 lbgidl = 344.995831 wbgidl = -3.677361E3
+ pbgidl = 7.021001E-3 cgidl = 78.73687 lcgidl = 7.442507E-4
+ wcgidl = 7.206757E-3 pcgidl = -1.37595E-8 egidl = 3.110213
+ legidl = -2.119675E-6 noia = 3E40 noib = 8.53E24
+ noic = 8.4E7 em = 4.1E7 af = 1
+ ef = 0.88 kf = 0 lintnoi = 0
+ tnoia = 1.5 tnoib = 3.5 ntnoi = 1
+ rnoia = 0.577 rnoib = 0.37 xpart = 0
+ cgso = {1.94171E-10/sw_func_tox_hv_ratio} cgdo = {1.94171E-10/sw_func_tox_hv_ratio} cgbo = {0/sw_func_tox_hv_ratio}
+ ckappas = 0.6 cf = 1.2E-11 clc = 1E-7
+ cle = 0.6 dlc = 4.4983E-8 dwc = 0
+ vfbcv = -0.144689 noff = 4 voffcv = 0
+ acde = 0.401 moin = 15.773 cgsl = {9.82591E-12/sw_func_tox_hv_ratio}
+ cgdl = {9.82591E-12/sw_func_tox_hv_ratio} ijthsrev = 0.1 ijthsfwd = 0.1
+ xjbvs = 1 bvs = 12.69 jss = 2.1483E-5
+ jsws = 4.02E-12 cjs = {sw_psd_nw_cj} mjs = 0.33956
+ mjsws = 0.24676 cjsws = {9.960545E-11*sw_func_psd_nw_cj} cjswgs = {1.47314E-10*sw_func_psd_nw_cj}
+ mjswgs = 0.81 pbs = 0.6587 pbsws = 1
+ pbswgs = 3 xrcrg1 = 12 xrcrg2 = 1
+ rbpb = 50 rbpd = 50 rbps = 50
+ rbdb = 50 rbsb = 50 gbmin = 1E-12
+ tnom = 30 ute = -1.211876 lute = -3.591754E-7
+ kt1 = -0.513878 lkt1 = -9.760501E-8 wkt1 = 2.719941E-7
+ pkt1 = -5.193048E-13 kt1l = 0 kt2 = -0.019032
+ ua1 = 6.729484E-10 lua1 = -2.30157E-16 ub1 = -3.532041E-18
+ lub1 = -2.494611E-25 uc1 = -1.092E-10 at = 2.662658E5
+ lat = -0.220453 wat = -0.108798 pat = 2.077219E-7
+ prt = 0 njs = 1.3632 xtis = 10
+ tpb = 1.671E-3 tpbsw = 0 tpbswg = 0
+ tcj = 9.6E-4 tcjsw = 3E-5 tcjswg = 0
+ tvoff = 0 tvfbsdoff = 0 saref = 3E-6
+ sbref = 3E-6 wlod = 0 ku0 = 7E-8
+ kvsat = 0.4 kvth0 = 3.5E-8 tku0 = 0
+ llodku0 = 0 wlodku0 = 1 llodvth = 0
+ wlodvth = 1 lku0 = 0 wku0 = 0
+ pku0 = 0 lkvth0 = 0 wkvth0 = 6.5E-7
+ pkvth0 = 0 stk2 = 0 lodk2 = 1
+ steta0 = 0 lodeta0 = 1

.model phv_model.12 pmos
+ level = 54 lmin = 8E-7 lmax = 1E-6 wmin = 1.5E-5
+ wmax = 2E-5 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 1.175E-8
+ toxm = 1.175E-8 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 1E23 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {1.2277E-8+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {4.5375E-8-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = -4.7338E-9 dwb = 0 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = -1.136948 lvth0 = 1.162593E-7
+ wvth0 = 1.007738E-6 pvth0 = -7.147384E-13 k1 = 0.590242
+ lk1 = -9.866749E-9 k2 = 2.03531E-2 lk2 = 1.132523E-8
+ wk2 = 3.753519E-8 pk2 = -2.662184E-14 k3 = -2.2405
+ k3b = -0.172 w0 = 0 lpe0 = 0
+ lpeb = 0 vbm = -3 dvtp0 = 0
+ dvtp1 = 0 dvt0 = 4.657 dvt1 = 0.34864
+ dvt2 = -0.030206 dvt0w = -2.2 dvt1w = 1.0163E6
+ dvt2w = 0 vfbsdoff = 0 u0 = 2.16928E-2
+ lu0 = -1.787576E-9 wu0 = -5.064531E-8 pu0 = 3.592019E-14
+ ua = -8.10062E-10 lua = 2.239702E-15 wua = -2.092206E-16
+ pua = 1.483897E-22 ub = 4.770673E-18 lub = -3.504144E-24
+ wub = -8.3611E-24 pub = 5.93011E-30 uc = 6.082696E-12
+ luc = -6.063021E-18 ud = 0 up = 0
+ lp = 1 eu = 1.67 vsat = 8.367108E3
+ lvsat = 3.59353E-2 a0 = 0.797865 la0 = 3.237399E-8
+ wa0 = -6.799854E-8 pa0 = 4.822796E-14 ags = 0.768933
+ lags = -3.391159E-8 wags = 3.924876E-7 pags = -2.783718E-13
+ b0 = 0 b1 = 0 keta = -0.15376
+ lketa = 6.28183E-8 a1 = 0 a2 = 0.5
+ rdsw = 788.47 rdswmin = 0 rdw = 0
+ rdwmin = 0 rsw = 0 rswmin = 0
+ prwb = 0.053538 prwg = 0 wr = 1
+ voff = -9.52546E-2 lvoff = 1.591078E-8 voffl = 0
+ minv = 0 nfactor = 0.77916 lnfactor = 6.335166E-7
+ wnfactor = 8.080946E-6 pnfactor = -5.731411E-12 eta0 = -2.551868E-4
+ leta0 = 2.21366E-10 weta0 = 3.665937E-9 peta0 = -2.600066E-15
+ etab = 7.545356E-4 letab = -6.860615E-10 dsub = 1.499307
+ ldsub = -8.684674E-7 cit = -1.273125E-5 lcit = 1.612214E-11
+ cdsc = 0 cdscb = 0 cdscd = 0
+ pclm = 2.021902 lpclm = -7.444957E-7 pdiblc1 = 0.195862
+ lpdiblc1 = 1.851818E-7 pdiblc2 = -3.36185E-2 lpdiblc2 = 3.193712E-8
+ pdiblcb = -0.025 drout = 0.335842 ldrout = 6.805458E-8
+ pscbe1 = -5.698769E7 lpscbe1 = 324.118516 pscbe2 = 1.828151E-8
+ lpscbe2 = -3.388725E-15 pvag = 0 delta = 0.01
+ fprout = 0 pdits = 0 pditsl = 0
+ pditsd = 0 lambda = 0 vtl = 0
+ lc = 5E-9 xn = 3 alpha0 = 2.471576E-4
+ lalpha0 = -1.63069E-10 alpha1 = 0 beta0 = 67.196894
+ lbeta0 = -1.549723E-5 aigbacc = 0.43 bigbacc = 0.054
+ cigbacc = 0.075 nigbacc = 1 aigbinv = 0.35
+ bigbinv = 0.03 cigbinv = 6E-3 eigbinv = 1.1
+ nigbinv = 3 aigc = 0.43 bigc = 0.054
+ cigc = 0.075 aigsd = 0.43 bigsd = 0.054
+ cigsd = 0.075 dlcig = 0 nigc = 1
+ poxedge = 1 pigcd = 1 ntox = 1
+ toxref = 1.175E-8 agidl = 4.313149E-8 lagidl = -2.253393E-14
+ wagidl = -6.809645E-13 pagidl = 4.829741E-19 bgidl = 4.122722E7
+ lbgidl = 1.252587E3 wbgidl = 1.83868E4 pbgidl = -1.30408E-2
+ cgidl = 2.235161E3 lcgidl = -1.216478E-3 wcgidl = -3.60338E-2
+ pcgidl = 2.555696E-8 egidl = 1.835557 legidl = -9.606931E-7
+ noia = 3E40 noib = 8.53E24 noic = 8.4E7
+ em = 4.1E7 af = 1 ef = 0.88
+ kf = 0 lintnoi = 0 tnoia = 1.5
+ tnoib = 3.5 ntnoi = 1 rnoia = 0.577
+ rnoib = 0.37 xpart = 0 cgso = {1.94171E-10/sw_func_tox_hv_ratio}
+ cgdo = {1.94171E-10/sw_func_tox_hv_ratio} cgbo = {0/sw_func_tox_hv_ratio} ckappas = 0.6
+ cf = 1.2E-11 clc = 1E-7 cle = 0.6
+ dlc = 4.4983E-8 dwc = 0 vfbcv = -0.144689
+ noff = 4 voffcv = 0 acde = 0.401
+ moin = 15.773 cgsl = {9.82591E-12/sw_func_tox_hv_ratio} cgdl = {9.82591E-12/sw_func_tox_hv_ratio}
+ ijthsrev = 0.1 ijthsfwd = 0.1 xjbvs = 1
+ bvs = 12.69 jss = 2.1483E-5 jsws = 4.02E-12
+ cjs = {sw_psd_nw_cj} mjs = 0.33956 mjsws = 0.24676
+ cjsws = {9.960545E-11*sw_func_psd_nw_cj} cjswgs = {1.47314E-10*sw_func_psd_nw_cj} mjswgs = 0.81
+ pbs = 0.6587 pbsws = 1 pbswgs = 3
+ xrcrg1 = 12 xrcrg2 = 1 rbpb = 50
+ rbpd = 50 rbps = 50 rbdb = 50
+ rbsb = 50 gbmin = 1E-12 tnom = 30
+ ute = -2.057628 lute = 4.098248E-7 kt1 = -0.54223
+ lkt1 = -7.182557E-8 wkt1 = -1.359971E-6 pkt1 = 9.645592E-13
+ kt1l = 0 kt2 = -0.019032 ua1 = -5.034182E-11
+ lua1 = 4.274946E-16 ub1 = -4.570617E-18 lub1 = 6.948642E-25
+ uc1 = -1.092E-10 at = 1.958915E4 lat = 3.837644E-3
+ wat = 0.543988 pat = -3.858237E-7 prt = 0
+ njs = 1.3632 xtis = 10 tpb = 1.671E-3
+ tpbsw = 0 tpbswg = 0 tcj = 9.6E-4
+ tcjsw = 3E-5 tcjswg = 0 tvoff = 0
+ tvfbsdoff = 0 saref = 2.81E-6 sbref = 2.81E-6
+ wlod = 0 ku0 = 7E-8 kvsat = 0.4
+ kvth0 = 3.5E-8 tku0 = 0 llodku0 = 0
+ wlodku0 = 1 llodvth = 0 wlodvth = 1
+ lku0 = 0 wku0 = 0 pku0 = 0
+ lkvth0 = 0 wkvth0 = 6.5E-7 pkvth0 = 0
+ stk2 = 0 lodk2 = 1 steta0 = 0
+ lodeta0 = 1

.model phv_model.13 pmos
+ level = 54 lmin = 6E-7 lmax = 8E-7 wmin = 1.5E-5
+ wmax = 2E-5 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 1.175E-8
+ toxm = 1.175E-8 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 1E23 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {1.2277E-8+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {4.5375E-8-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = -4.7338E-9 dwb = 0 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = -0.973029 k1 = 0.57633
+ k2 = 0.036321 k3 = -2.2405 k3b = -0.172
+ w0 = 0 lpe0 = 0 lpeb = 0
+ vbm = -3 dvtp0 = 0 dvtp1 = 0
+ dvt0 = 4.657 dvt1 = 0.34864 dvt2 = -0.030206
+ dvt0w = -2.2 dvt1w = 1.0163E6 dvt2w = 0
+ vfbsdoff = 0 u0 = 1.91724E-2 ua = 2.347784E-9
+ ub = -1.6996E-19 uc = -2.4658E-12 ud = 0
+ up = 0 lp = 1 eu = 1.67
+ vsat = 5.90337E4 a0 = 0.84351 ags = 0.72112
+ b0 = 0 b1 = 0 keta = -0.06519
+ a1 = 0 a2 = 0.5 rdsw = 788.47
+ rdswmin = 0 rdw = 0 rdwmin = 0
+ rsw = 0 rswmin = 0 prwb = 0.053538
+ prwg = 0 wr = 1 voff = -7.28213E-2
+ voffl = 0 minv = 0 nfactor = 1.67238
+ eta0 = 5.6926E-5 etab = -2.1277E-4 dsub = 0.27482
+ cit = 1E-5 cdsc = 0 cdscb = 0
+ cdscd = 0 pclm = 0.972208 pdiblc1 = 0.456957
+ pdiblc2 = 1.14109E-2 pdiblcb = -0.025 drout = 0.431795
+ pscbe1 = 4E8 pscbe2 = 1.350362E-8 pvag = 0
+ delta = 0.01 fprout = 0 pdits = 0
+ pditsl = 0 pditsd = 0 lambda = 0
+ vtl = 0 lc = 5E-9 xn = 3
+ alpha0 = 1.724017E-5 alpha1 = 0 beta0 = 45.34673
+ aigbacc = 0.43 bigbacc = 0.054 cigbacc = 0.075
+ nigbacc = 1 aigbinv = 0.35 bigbinv = 0.03
+ cigbinv = 6E-3 eigbinv = 1.1 nigbinv = 3
+ aigc = 0.43 bigc = 0.054 cigc = 0.075
+ aigsd = 0.43 bigsd = 0.054 cigsd = 0.075
+ dlcig = 0 nigc = 1 poxedge = 1
+ pigcd = 1 ntox = 1 toxref = 1.175E-8
+ agidl = 1.136E-8 bgidl = 1.8073E9 cgidl = 520
+ egidl = 0.481037 noia = 3E40 noib = 8.53E24
+ noic = 8.4E7 em = 4.1E7 af = 1
+ ef = 0.88 kf = 0 lintnoi = 0
+ tnoia = 1.5 tnoib = 3.5 ntnoi = 1
+ rnoia = 0.577 rnoib = 0.37 xpart = 0
+ cgso = {1.94171E-10/sw_func_tox_hv_ratio} cgdo = {1.94171E-10/sw_func_tox_hv_ratio} cgbo = {0/sw_func_tox_hv_ratio}
+ ckappas = 0.6 cf = 1.2E-11 clc = 1E-7
+ cle = 0.6 dlc = 4.4983E-8 dwc = 0
+ vfbcv = -0.144689 noff = 4 voffcv = 0
+ acde = 0.401 moin = 15.773 cgsl = {9.82591E-12/sw_func_tox_hv_ratio}
+ cgdl = {9.82591E-12/sw_func_tox_hv_ratio} ijthsrev = 0.1 ijthsfwd = 0.1
+ xjbvs = 1 bvs = 12.69 jss = 2.1483E-5
+ jsws = 4.02E-12 cjs = {sw_psd_nw_cj} mjs = 0.33956
+ mjsws = 0.24676 cjsws = {9.960545E-11*sw_func_psd_nw_cj} cjswgs = {1.47314E-10*sw_func_psd_nw_cj}
+ mjswgs = 0.81 pbs = 0.6587 pbsws = 1
+ pbswgs = 3 xrcrg1 = 12 xrcrg2 = 1
+ rbpb = 50 rbpd = 50 rbps = 50
+ rbdb = 50 rbsb = 50 gbmin = 1E-12
+ tnom = 30 ute = -1.4798 kt1 = -0.6435
+ kt1l = 0 kt2 = -0.019032 ua1 = 5.524E-10
+ ub1 = -3.5909E-18 uc1 = -1.092E-10 at = 2.5E4
+ prt = 0 njs = 1.3632 xtis = 10
+ tpb = 1.671E-3 tpbsw = 0 tpbswg = 0
+ tcj = 9.6E-4 tcjsw = 3E-5 tcjswg = 0
+ tvoff = 0 tvfbsdoff = 0 saref = 2.41E-6
+ sbref = 2.41E-6 wlod = 0 ku0 = 7E-8
+ kvsat = 0.4 kvth0 = 3.5E-8 tku0 = 0
+ llodku0 = 0 wlodku0 = 1 llodvth = 0
+ wlodvth = 1 lku0 = 0 wku0 = 0
+ pku0 = 0 lkvth0 = 0 wkvth0 = 6.5E-7
+ pkvth0 = 0 stk2 = 0 lodk2 = 1
+ steta0 = 0 lodeta0 = 1

.model phv_model.14 pmos
+ level = 54 lmin = 5E-7 lmax = 6E-7 wmin = 1.5E-5
+ wmax = 2E-5 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 1.175E-8
+ toxm = 1.175E-8 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 1E23 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {1.2277E-8+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {4.5375E-8-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = -4.7338E-9 dwb = 0 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = -0.739554 lvth0 = -1.188972E-7
+ wvth0 = -8.731247E-7 pvth0 = 4.446388E-13 k1 = 0.487482
+ lk1 = 4.524593E-8 k2 = 2.70453E-2 lk2 = 4.723654E-9
+ wk2 = 2.423986E-8 pk2 = -1.234415E-14 k3 = -2.2405
+ k3b = -0.172 w0 = 0 lpe0 = 0
+ lpeb = 0 vbm = -3 dvtp0 = 0
+ dvtp1 = 0 dvt0 = 4.657 dvt1 = 0.34864
+ dvt2 = -0.030206 dvt0w = -2.2 dvt1w = 1.0163E6
+ dvt2w = 0 vfbsdoff = 0 u0 = 0.010551
+ lu0 = 4.390471E-9 wu0 = 5.259315E-8 pu0 = -2.678306E-14
+ ua = 3.107579E-9 lua = -3.869259E-16 wua = 1.669147E-16
+ pua = -8.500131E-23 ub = -3.145609E-18 lub = 1.515349E-24
+ wub = -1.897565E-24 pub = 9.663349E-31 uc = 9.057452E-12
+ luc = -5.868216E-18 ud = 0 up = 0
+ lp = 1 eu = 1.67 vsat = 4.861593E4
+ lvsat = 5.305248E-3 wvsat = -0.113438 pvsat = 5.776813E-8
+ a0 = 0.368248 la0 = 2.420272E-7 ags = -1.443321
+ lags = 1.102242E-6 b0 = 0 b1 = 0
+ keta = 1.94429E-2 lketa = -4.30993E-8 a1 = 0
+ a2 = 0.5 rdsw = 788.47 rdswmin = 0
+ rdw = 0 rdwmin = 0 rsw = 0
+ rswmin = 0 prwb = 0.053538 prwg = 0
+ wr = 1 voff = 4.46966E-2 lvoff = -5.984601E-8
+ voffl = 0 minv = 0 nfactor = 2.104033
+ lnfactor = -2.198195E-7 wnfactor = -8.263589E-6 pnfactor = 4.208233E-12
+ eta0 = -0.464716 leta0 = 2.366857E-7 weta0 = 2.744246E-6
+ peta0 = -1.397507E-12 etab = 1.46738E-2 letab = -7.580997E-9
+ dsub = 0.254971 ldsub = 1.010791E-8 cit = 3.04625E-5
+ lcit = -1.042053E-11 cdsc = 0 cdscb = 0
+ cdscd = 0 pclm = -0.519068 lpclm = 7.594321E-7
+ pdiblc1 = 1.123736 lpdiblc1 = -3.39557E-7 pdiblc2 = 3.84625E-2
+ lpdiblc2 = -1.377603E-8 pdiblcb = -0.025 drout = -1.482714
+ ldrout = 9.749638E-7 pscbe1 = 5.52896E8 lpscbe1 = -77.86227
+ pscbe2 = 9.480217E-9 lpscbe2 = 2.048916E-15 pvag = 0
+ delta = 0.01 fprout = 0 pdits = 0
+ pditsl = 0 pditsd = 0 lambda = 0
+ vtl = 0 lc = 5E-9 xn = 3
+ alpha0 = -3.097308E-4 lalpha0 = 1.6651E-10 alpha1 = 0
+ beta0 = 7.131861 lbeta0 = 1.946092E-5 aigbacc = 0.43
+ bigbacc = 0.054 cigbacc = 0.075 nigbacc = 1
+ aigbinv = 0.35 bigbinv = 0.03 cigbinv = 6E-3
+ eigbinv = 1.1 nigbinv = 3 aigc = 0.43
+ bigc = 0.054 cigc = 0.075 aigsd = 0.43
+ bigsd = 0.054 cigsd = 0.075 dlcig = 0
+ nigc = 1 poxedge = 1 pigcd = 1
+ ntox = 1 toxref = 1.175E-8 agidl = -1.682469E-9
+ lagidl = 6.641877E-15 wagidl = 5.386636E-14 pagidl = -2.743144E-20
+ bgidl = 2.657621E9 lbgidl = -433.025976 wbgidl = -1.224235E3
+ pbgidl = 6.234419E-4 cgidl = -7.79274E3 lcgidl = 4.233263E-3
+ wcgidl = 0.136948 pcgidl = -6.97407E-8 egidl = -0.272932
+ legidl = 3.839585E-7 noia = 3E40 noib = 8.53E24
+ noic = 8.4E7 em = 4.1E7 af = 1
+ ef = 0.88 kf = 0 lintnoi = 0
+ tnoia = 1.5 tnoib = 3.5 ntnoi = 1
+ rnoia = 0.577 rnoib = 0.37 xpart = 0
+ cgso = {1.94171E-10/sw_func_tox_hv_ratio} cgdo = {1.94171E-10/sw_func_tox_hv_ratio} cgbo = {0/sw_func_tox_hv_ratio}
+ ckappas = 0.6 cf = 1.2E-11 clc = 1E-7
+ cle = 0.6 dlc = 4.4983E-8 dwc = 0
+ vfbcv = -0.144689 noff = 4 voffcv = 0
+ acde = 0.401 moin = 15.773 cgsl = {9.82591E-12/sw_func_tox_hv_ratio}
+ cgdl = {9.82591E-12/sw_func_tox_hv_ratio} ijthsrev = 0.1 ijthsfwd = 0.1
+ xjbvs = 1 bvs = 12.69 jss = 2.1483E-5
+ jsws = 4.02E-12 cjs = {sw_psd_nw_cj} mjs = 0.33956
+ mjsws = 0.24676 cjsws = {9.960545E-11*sw_func_psd_nw_cj} cjswgs = {1.47314E-10*sw_func_psd_nw_cj}
+ mjswgs = 0.81 pbs = 0.6587 pbsws = 1
+ pbswgs = 3 xrcrg1 = 12 xrcrg2 = 1
+ rbpb = 50 rbpd = 50 rbps = 50
+ rbdb = 50 rbsb = 50 gbmin = 1E-12
+ tnom = 30 ute = -1.919334 lute = 2.238329E-7
+ kt1 = -0.643783 lkt1 = 1.440284E-10 wkt1 = -2.448471E-6
+ pkt1 = 1.246884E-12 kt1l = 0 kt2 = -0.019032
+ ua1 = 5.524E-10 ub1 = -9.446858E-18 lub1 = 2.982147E-24
+ uc1 = -3.862786E-10 luc1 = 1.411023E-16 at = 5.36475E4
+ lat = -1.45887E-2 prt = 0 njs = 1.3632
+ xtis = 10 tpb = 1.671E-3 tpbsw = 0
+ tpbswg = 0 tcj = 9.6E-4 tcjsw = 3E-5
+ tcjswg = 0 tvoff = 0 tvfbsdoff = 0
+ saref = 2.41E-6 sbref = 2.41E-6 wlod = 0
+ ku0 = 7E-8 kvsat = 0.4 kvth0 = 3.5E-8
+ tku0 = 0 llodku0 = 0 wlodku0 = 1
+ llodvth = 0 wlodvth = 1 lku0 = 0
+ wku0 = 0 pku0 = 0 lkvth0 = 0
+ wkvth0 = 6.5E-7 pkvth0 = 0 stk2 = 0
+ lodk2 = 1 steta0 = 0 lodeta0 = 1

.model phv_model.15 pmos
+ level = 54 lmin = 8E-6 lmax = 2.02E-5 wmin = 7E-6
+ wmax = 1.5E-5 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 1.175E-8
+ toxm = 1.175E-8 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 1E23 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {1.2277E-8+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {4.5375E-8-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = -4.7338E-9 dwb = 0 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = -1.011028 k1 = 0.59521
+ k2 = 2.52804E-2 k3 = -2.2405 k3b = -0.172
+ w0 = 0 lpe0 = 0 lpeb = 0
+ vbm = -3 dvtp0 = 0 dvtp1 = 0
+ dvt0 = 4.657 dvt1 = 0.34864 dvt2 = -0.030206
+ dvt0w = -2.2 dvt1w = 1.0163E6 dvt2w = 0
+ vfbsdoff = 0 u0 = 2.09856E-2 ua = 2.704411E-9
+ ub = -1.7524E-19 uc = -3.9972E-11 ud = 0
+ up = 0 lp = 1 eu = 1.67
+ vsat = 2E5 a0 = 0.89674 ags = 0.134273
+ b0 = 0 b1 = 0 keta = -7.9259E-3
+ a1 = 0 a2 = 0.5 rdsw = 788.47
+ rdswmin = 0 rdw = 0 rdwmin = 0
+ rsw = 0 rswmin = 0 prwb = 0.053538
+ prwg = 0 wr = 1 voff = -9.32047E-2
+ voffl = 0 minv = 0 nfactor = 1.74009
+ eta0 = 0.08 etab = -0.07 dsub = 0.56
+ cit = 1E-5 cdsc = 0 cdscb = 0
+ cdscd = 0 pclm = 8.35312E-2 pdiblc1 = 0.39
+ pdiblc2 = 2.940788E-3 pdiblcb = -0.025 drout = 0.56
+ pscbe1 = 3.337128E8 pscbe2 = 1.500096E-8 pvag = 0
+ delta = 0.01 fprout = 0 pdits = 0
+ pditsl = 0 pditsd = 0 lambda = 0
+ vtl = 0 lc = 5E-9 xn = 3
+ alpha0 = 5.066719E-5 alpha1 = 0 beta0 = 38.266046
+ aigbacc = 0.43 bigbacc = 0.054 cigbacc = 0.075
+ nigbacc = 1 aigbinv = 0.35 bigbinv = 0.03
+ cigbinv = 6E-3 eigbinv = 1.1 nigbinv = 3
+ aigc = 0.43 bigc = 0.054 cigc = 0.075
+ aigsd = 0.43 bigsd = 0.054 cigsd = 0.075
+ dlcig = 0 nigc = 1 poxedge = 1
+ pigcd = 1 ntox = 1 toxref = 1.175E-8
+ agidl = 7.3657E-9 bgidl = 1.7047E9 cgidl = 700
+ egidl = 0.693508 noia = 3E40 noib = 8.53E24
+ noic = 8.4E7 em = 4.1E7 af = 1
+ ef = 0.88 kf = 0 lintnoi = 0
+ tnoia = 1.5 tnoib = 3.5 ntnoi = 1
+ rnoia = 0.577 rnoib = 0.37 xpart = 0
+ cgso = {1.94171E-10/sw_func_tox_hv_ratio} cgdo = {1.94171E-10/sw_func_tox_hv_ratio} cgbo = {0/sw_func_tox_hv_ratio}
+ ckappas = 0.6 cf = 1.2E-11 clc = 1E-7
+ cle = 0.6 dlc = 4.4983E-8 dwc = 0
+ vfbcv = -0.144689 noff = 4 voffcv = 0
+ acde = 0.401 moin = 15.773 cgsl = {9.82591E-12/sw_func_tox_hv_ratio}
+ cgdl = {9.82591E-12/sw_func_tox_hv_ratio} ijthsrev = 0.1 ijthsfwd = 0.1
+ xjbvs = 1 bvs = 12.69 jss = 2.1483E-5
+ jsws = 4.02E-12 cjs = {sw_psd_nw_cj} mjs = 0.33956
+ mjsws = 0.24676 cjsws = {9.960545E-11*sw_func_psd_nw_cj} cjswgs = {1.47314E-10*sw_func_psd_nw_cj}
+ mjswgs = 0.81 pbs = 0.6587 pbsws = 1
+ pbswgs = 3 xrcrg1 = 12 xrcrg2 = 1
+ rbpb = 50 rbpd = 50 rbps = 50
+ rbdb = 50 rbsb = 50 gbmin = 1E-12
+ tnom = 30 ute = -1.3864 kt1 = -0.57573
+ kt1l = 0 kt2 = -0.019032 ua1 = 7.0656E-10
+ ub1 = -3.145E-18 uc1 = -1.092E-10 at = 4.3E5
+ prt = 0 njs = 1.3632 xtis = 10
+ tpb = 1.671E-3 tpbsw = 0 tpbswg = 0
+ tcj = 9.6E-4 tcjsw = 3E-5 tcjswg = 0
+ tvoff = 0 tvfbsdoff = 0 saref = 3E-6
+ sbref = 3E-6 wlod = 0 ku0 = 7E-8
+ kvsat = 0.4 kvth0 = 3.5E-8 tku0 = 0
+ llodku0 = 0 wlodku0 = 1 llodvth = 0
+ wlodvth = 1 lku0 = 0 wku0 = 0
+ pku0 = 0 lkvth0 = 0 wkvth0 = 6.5E-7
+ pkvth0 = 0 stk2 = 0 lodk2 = 1
+ steta0 = 0 lodeta0 = 1

.model phv_model.16 pmos
+ level = 54 lmin = 4E-6 lmax = 8E-6 wmin = 7E-6
+ wmax = 1.5E-5 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 1.175E-8
+ toxm = 1.175E-8 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 1E23 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {1.2277E-8+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {4.5375E-8-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = -4.7338E-9 dwb = 0 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = -1.016266 lvth0 = 4.143178E-8
+ k1 = 0.604152 lk1 = -7.072775E-8 k2 = 2.32995E-2
+ lk2 = 1.566755E-8 k3 = -2.2405 k3b = -0.172
+ w0 = 0 lpe0 = 0 lpeb = 0
+ vbm = -3 dvtp0 = 0 dvtp1 = 0
+ dvt0 = 4.657 dvt1 = 0.34864 dvt2 = -0.030206
+ dvt0w = -2.2 dvt1w = 1.0163E6 dvt2w = 0
+ vfbsdoff = 0 u0 = 2.02516E-2 lu0 = 5.805086E-9
+ ua = 2.449766E-9 lua = 2.014057E-15 ub = 8.85171E-20
+ lub = -2.086121E-24 uc = -5.157563E-11 luc = 9.177602E-17
+ ud = 0 up = 0 lp = 1
+ eu = 1.67 vsat = 2.977215E5 lvsat = -0.772904
+ a0 = 0.916542 la0 = -1.566198E-7 ags = 0.109759
+ lags = 1.93893E-7 b0 = 0 b1 = 0
+ keta = -4.956727E-3 lketa = -2.348393E-8 a1 = 0
+ a2 = 0.5 rdsw = 788.47 rdswmin = 0
+ rdw = 0 rdwmin = 0 rsw = 0
+ rswmin = 0 prwb = 0.053538 prwg = 0
+ wr = 1 voff = -9.47765E-2 lvoff = 1.243193E-8
+ voffl = 0 minv = 0 nfactor = 1.75518
+ lnfactor = -1.193482E-7 eta0 = 0.08 etab = -0.07
+ dsub = 0.56 cit = 1E-5 cdsc = 0
+ cdscb = 0 cdscd = 0 pclm = -0.648319
+ lpclm = 5.788389E-6 pdiblc1 = 0.39 pdiblc2 = 4.554123E-3
+ lpdiblc2 = -1.276027E-8 pdiblcb = -0.025 drout = 0.56
+ pscbe1 = 5.621233E8 lpscbe1 = -1.806556E3 pscbe2 = -1.531739E-8
+ lpscbe2 = 2.397954E-13 pvag = 0 delta = 0.01
+ fprout = 0 pdits = 0 pditsl = 0
+ pditsd = 0 lambda = 0 vtl = 0
+ lc = 5E-9 xn = 3 alpha0 = 7.815322E-5
+ lalpha0 = -2.173939E-10 alpha1 = 0 beta0 = 39.140288
+ lbeta0 = -6.9146E-6 aigbacc = 0.43 bigbacc = 0.054
+ cigbacc = 0.075 nigbacc = 1 aigbinv = 0.35
+ bigbinv = 0.03 cigbinv = 6E-3 eigbinv = 1.1
+ nigbinv = 3 aigc = 0.43 bigc = 0.054
+ cigc = 0.075 aigsd = 0.43 bigsd = 0.054
+ cigsd = 0.075 dlcig = 0 nigc = 1
+ poxedge = 1 pigcd = 1 ntox = 1
+ toxref = 1.175E-8 agidl = 6.538796E-9 lagidl = 6.540191E-15
+ bgidl = 1.478354E9 lbgidl = 1.790224E3 cgidl = 932.600375
+ lcgidl = -1.839695E-3 egidl = 1.209319 legidl = -4.079675E-6
+ noia = 3E40 noib = 8.53E24 noic = 8.4E7
+ em = 4.1E7 af = 1 ef = 0.88
+ kf = 0 lintnoi = 0 tnoia = 1.5
+ tnoib = 3.5 ntnoi = 1 rnoia = 0.577
+ rnoib = 0.37 xpart = 0 cgso = {1.94171E-10/sw_func_tox_hv_ratio}
+ cgdo = {1.94171E-10/sw_func_tox_hv_ratio} cgbo = {0/sw_func_tox_hv_ratio} ckappas = 0.6
+ cf = 1.2E-11 clc = 1E-7 cle = 0.6
+ dlc = 4.4983E-8 dwc = 0 vfbcv = -0.144689
+ noff = 4 voffcv = 0 acde = 0.401
+ moin = 15.773 cgsl = {9.82591E-12/sw_func_tox_hv_ratio} cgdl = {9.82591E-12/sw_func_tox_hv_ratio}
+ ijthsrev = 0.1 ijthsfwd = 0.1 xjbvs = 1
+ bvs = 12.69 jss = 2.1483E-5 jsws = 4.02E-12
+ cjs = {sw_psd_nw_cj} mjs = 0.33956 mjsws = 0.24676
+ cjsws = {9.960545E-11*sw_func_psd_nw_cj} cjswgs = {1.47314E-10*sw_func_psd_nw_cj} mjswgs = 0.81
+ pbs = 0.6587 pbsws = 1 pbswgs = 3
+ xrcrg1 = 12 xrcrg2 = 1 rbpb = 50
+ rbpd = 50 rbps = 50 rbdb = 50
+ rbsb = 50 gbmin = 1E-12 tnom = 30
+ ute = -1.22055 lute = -1.311749E-6 kt1 = -0.585239
+ lkt1 = 7.521104E-8 kt1l = 0 kt2 = -0.019032
+ ua1 = 1.375495E-9 lua1 = -5.290776E-15 ub1 = -2.61041E-18
+ lub1 = -4.228205E-24 uc1 = -1.092E-10 at = 6.730478E5
+ lat = -1.922326 prt = 0 njs = 1.3632
+ xtis = 10 tpb = 1.671E-3 tpbsw = 0
+ tpbswg = 0 tcj = 9.6E-4 tcjsw = 3E-5
+ tcjswg = 0 tvoff = 0 tvfbsdoff = 0
+ saref = 3E-6 sbref = 3E-6 wlod = 0
+ ku0 = 7E-8 kvsat = 0.4 kvth0 = 3.5E-8
+ tku0 = 0 llodku0 = 0 wlodku0 = 1
+ llodvth = 0 wlodvth = 1 lku0 = 0
+ wku0 = 0 pku0 = 0 lkvth0 = 0
+ wkvth0 = 6.5E-7 pkvth0 = 0 stk2 = 0
+ lodk2 = 1 steta0 = 0 lodeta0 = 1

.model phv_model.17 pmos
+ level = 54 lmin = 2E-6 lmax = 4E-6 wmin = 7E-6
+ wmax = 1.5E-5 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 1.175E-8
+ toxm = 1.175E-8 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 1E23 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {1.2277E-8+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {4.5375E-8-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = -4.7338E-9 dwb = 0 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = -0.991137 lvth0 = -5.680649E-8
+ k1 = 0.602594 lk1 = -6.463595E-8 k2 = 2.68321E-2
+ lk2 = 1.857724E-9 k3 = -2.2405 k3b = -0.172
+ w0 = 0 lpe0 = 0 lpeb = 0
+ vbm = -3 dvtp0 = 0 dvtp1 = 0
+ dvt0 = 4.657 dvt1 = 0.34864 dvt2 = -0.030206
+ dvt0w = -2.2 dvt1w = 1.0163E6 dvt2w = 0
+ vfbsdoff = 0 u0 = 2.09383E-2 lu0 = 3.120588E-9
+ ua = 3.313866E-9 lua = -1.363927E-15 ub = -1.459991E-18
+ lub = 3.967386E-24 uc = -5.492301E-11 luc = 1.048618E-16
+ ud = 0 up = 0 lp = 1
+ eu = 1.67 vsat = 8.454508E4 lvsat = 6.04563E-2
+ a0 = 0.823723 la0 = 2.062331E-7 ags = 0.121307
+ lags = 1.487485E-7 b0 = 0 b1 = 0
+ keta = -5.087328E-3 lketa = -2.297338E-8 a1 = 0
+ a2 = 0.5 rdsw = 788.47 rdswmin = 0
+ rdw = 0 rdwmin = 0 rsw = 0
+ rswmin = 0 prwb = 0.053538 prwg = 0
+ wr = 1 voff = -0.064087 lvoff = -1.075408E-7
+ voffl = 0 minv = 0 nfactor = 2.156069
+ lnfactor = -1.686524E-6 eta0 = 1.90949E-2 leta0 = 2.380932E-7
+ etab = -0.122401 letab = 2.048497E-7 dsub = 0.814742
+ ldsub = -9.958489E-7 cit = 1E-5 cdsc = 0
+ cdscb = 0 cdscd = 0 pclm = 1.048766
+ lpclm = -8.459407E-7 pdiblc1 = 0.581562 lpdiblc1 = -7.488642E-7
+ pdiblc2 = -1.133342E-3 lpdiblc2 = 9.473451E-9 pdiblcb = 0.165925
+ lpdiblcb = -7.463736E-7 drout = 0.139965 ldrout = 1.642022E-6
+ pscbe1 = -1.561704E8 lpscbe1 = 1.001434E3 pscbe2 = 7.607469E-8
+ lpscbe2 = -1.174791E-13 pvag = 0 delta = 0.01
+ fprout = 0 pdits = 0 pditsl = 0
+ pditsd = 0 lambda = 0 vtl = 0
+ lc = 5E-9 xn = 3 alpha0 = 4.406319E-5
+ lalpha0 = -8.412745E-11 alpha1 = -9.54625E-11 lalpha1 = 3.731868E-16
+ beta0 = 70.183411 lbeta0 = -1.282699E-4 aigbacc = 0.43
+ bigbacc = 0.054 cigbacc = 0.075 nigbacc = 1
+ aigbinv = 0.35 bigbinv = 0.03 cigbinv = 6E-3
+ eigbinv = 1.1 nigbinv = 3 aigc = 0.43
+ bigc = 0.054 cigc = 0.075 aigsd = 0.43
+ bigsd = 0.054 cigsd = 0.075 dlcig = 0
+ nigc = 1 poxedge = 1 pigcd = 1
+ ntox = 1 toxref = 1.175E-8 agidl = 9.197164E-9
+ lagidl = -3.852034E-15 bgidl = 2.620002E9 lbgidl = -2.672764E3
+ cgidl = 455.747206 lcgidl = 2.444373E-5 egidl = -1.585323
+ legidl = 6.845277E-6 noia = 3E40 noib = 8.53E24
+ noic = 8.4E7 em = 4.1E7 af = 1
+ ef = 0.88 kf = 0 lintnoi = 0
+ tnoia = 1.5 tnoib = 3.5 ntnoi = 1
+ rnoia = 0.577 rnoib = 0.37 xpart = 0
+ cgso = {1.94171E-10/sw_func_tox_hv_ratio} cgdo = {1.94171E-10/sw_func_tox_hv_ratio} cgbo = {0/sw_func_tox_hv_ratio}
+ ckappas = 0.6 cf = 1.2E-11 clc = 1E-7
+ cle = 0.6 dlc = 4.4983E-8 dwc = 0
+ vfbcv = -0.144689 noff = 4 voffcv = 0
+ acde = 0.401 moin = 15.773 cgsl = {9.82591E-12/sw_func_tox_hv_ratio}
+ cgdl = {9.82591E-12/sw_func_tox_hv_ratio} ijthsrev = 0.1 ijthsfwd = 0.1
+ xjbvs = 1 bvs = 12.69 jss = 2.1483E-5
+ jsws = 4.02E-12 cjs = {sw_psd_nw_cj} mjs = 0.33956
+ mjsws = 0.24676 cjsws = {9.960545E-11*sw_func_psd_nw_cj} cjswgs = {1.47314E-10*sw_func_psd_nw_cj}
+ mjswgs = 0.81 pbs = 0.6587 pbsws = 1
+ pbswgs = 3 xrcrg1 = 12 xrcrg2 = 1
+ rbpb = 50 rbpd = 50 rbps = 50
+ rbdb = 50 rbsb = 50 gbmin = 1E-12
+ tnom = 30 ute = -1.705117 lute = 5.825446E-7
+ kt1 = -0.566955 lkt1 = 3.731868E-9 kt1l = 0
+ kt2 = -0.019032 ua1 = -4.841455E-10 lua1 = 1.979024E-15
+ ub1 = -3.719971E-18 lub1 = 1.093437E-25 uc1 = -1.092E-10
+ at = 2.104356E5 lat = -0.113859 prt = 0
+ njs = 1.3632 xtis = 10 tpb = 1.671E-3
+ tpbsw = 0 tpbswg = 0 tcj = 9.6E-4
+ tcjsw = 3E-5 tcjswg = 0 tvoff = 0
+ tvfbsdoff = 0 saref = 3E-6 sbref = 3E-6
+ wlod = 0 ku0 = 7E-8 kvsat = 0.4
+ kvth0 = 3.5E-8 tku0 = 0 llodku0 = 0
+ wlodku0 = 1 llodvth = 0 wlodvth = 1
+ lku0 = 0 wku0 = 0 pku0 = 0
+ lkvth0 = 0 wkvth0 = 6.5E-7 pkvth0 = 0
+ stk2 = 0 lodk2 = 1 steta0 = 0
+ lodeta0 = 1

.model phv_model.18 pmos
+ level = 54 lmin = 1E-6 lmax = 2E-6 wmin = 7E-6
+ wmax = 1.5E-5 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 1.175E-8
+ toxm = 1.175E-8 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 1E23 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {1.2277E-8+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {4.5375E-8-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = -4.7338E-9 dwb = 0 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = -1.034116 lvth0 = 2.525243E-8
+ wvth0 = -1.642215E-7 pvth0 = 3.135399E-13 k1 = 0.559056
+ lk1 = 1.848825E-8 k2 = 0.02248 lk2 = 1.016695E-8
+ wk2 = 4.107912E-9 pk2 = -7.843032E-15 k3 = -2.2405
+ k3b = -0.172 w0 = 0 lpe0 = 0
+ lpeb = 0 vbm = -3 dvtp0 = 0
+ dvtp1 = 0 dvt0 = 4.657 dvt1 = 0.34864
+ dvt2 = -0.030206 dvt0w = -2.2 dvt1w = 1.0163E6
+ dvt2w = 0 vfbsdoff = 0 u0 = 2.51653E-2
+ lu0 = -4.949794E-9 wu0 = 1.005726E-8 pu0 = -1.920183E-14
+ ua = 3.462173E-9 lua = -1.647083E-15 wua = 8.071141E-18
+ pua = -1.540983E-23 ub = 3.759318E-19 lub = 4.621496E-25
+ wub = 1.228574E-24 pub = -2.345656E-30 uc = 5.323295E-13
+ luc = -1.01635E-18 ud = 0 up = 0
+ lp = 1 eu = 1.67 vsat = 1.783309E5
+ lvsat = -0.118604 a0 = 1.01579 la0 = -1.604722E-7
+ wa0 = 9.300978E-8 pa0 = -1.775789E-13 ags = -0.299378
+ lags = 9.519411E-7 wags = 1.385055E-7 pags = -2.644416E-13
+ b0 = 0 b1 = 0 keta = 4.43017E-2
+ lketa = -1.172693E-7 a1 = 0 a2 = 0.5
+ rdsw = 788.47 rdswmin = 0 rdw = 0
+ rdwmin = 0 rsw = 0 rswmin = 0
+ prwb = 0.053538 prwg = 0 wr = 1
+ voff = -0.1592 lvoff = 7.405273E-8 voffl = 0
+ minv = 0 nfactor = 1.040892 lnfactor = 4.426273E-7
+ wnfactor = -9.10983E-7 pnfactor = 1.739294E-12 eta0 = 0.274512
+ leta0 = -2.495616E-7 etab = -2.88449E-2 letab = 2.622727E-8
+ dsub = 6.49192E-2 ldsub = 4.357497E-7 cit = 1.454625E-5
+ lcit = -8.679928E-12 cdsc = 0 cdscb = 0
+ cdscd = 0 pclm = 6.25064E-2 lpclm = 1.037075E-6
+ wpclm = -1.484072E-10 ppclm = 2.833465E-16 pdiblc1 = -1.786113E-3
+ lpdiblc1 = 3.648934E-7 pdiblc2 = 5.940119E-3 lpdiblc2 = -4.031554E-9
+ pdiblcb = -0.40685 lpdiblcb = 3.471971E-7 drout = 1.535831
+ ldrout = -1.023035E-6 pscbe1 = 4.309632E8 lpscbe1 = -119.550868
+ pscbe2 = 1.454314E-8 pvag = 0 delta = 0.01
+ fprout = 0 pdits = 0 pditsl = 0
+ pditsd = 0 lambda = 0 vtl = 0
+ lc = 5E-9 xn = 3 alpha0 = -6.165893E-5
+ lalpha0 = 1.177225E-10 alpha1 = 1.90925E-10 lalpha1 = -1.735986E-16
+ beta0 = -39.873797 lbeta0 = 8.18568E-5 aigbacc = 0.43
+ bigbacc = 0.054 cigbacc = 0.075 nigbacc = 1
+ aigbinv = 0.35 bigbinv = 0.03 cigbinv = 6E-3
+ eigbinv = 1.1 nigbinv = 3 aigc = 0.43
+ bigc = 0.054 cigc = 0.075 aigsd = 0.43
+ bigsd = 0.054 cigsd = 0.075 dlcig = 0
+ nigc = 1 poxedge = 1 pigcd = 1
+ ntox = 1 toxref = 1.175E-8 agidl = 6.118687E-9
+ lagidl = 2.025548E-15 bgidl = 7.938436E8 lbgidl = 813.830032
+ cgidl = 559.975088 lcgidl = -1.745533E-4 egidl = 3.110213
+ legidl = -2.119675E-6 noia = 3E40 noib = 8.53E24
+ noic = 8.4E7 em = 4.1E7 af = 1
+ ef = 0.88 kf = 0 lintnoi = 0
+ tnoia = 1.5 tnoib = 3.5 ntnoi = 1
+ rnoia = 0.577 rnoib = 0.37 xpart = 0
+ cgso = {1.94171E-10/sw_func_tox_hv_ratio} cgdo = {1.94171E-10/sw_func_tox_hv_ratio} cgbo = {0/sw_func_tox_hv_ratio}
+ ckappas = 0.6 cf = 1.2E-11 clc = 1E-7
+ cle = 0.6 dlc = 4.4983E-8 dwc = 0
+ vfbcv = -0.144689 noff = 4 voffcv = 0
+ acde = 0.401 moin = 15.773 cgsl = {9.82591E-12/sw_func_tox_hv_ratio}
+ cgdl = {9.82591E-12/sw_func_tox_hv_ratio} ijthsrev = 0.1 ijthsfwd = 0.1
+ xjbvs = 1 bvs = 12.69 jss = 2.1483E-5
+ jsws = 4.02E-12 cjs = {sw_psd_nw_cj} mjs = 0.33956
+ mjsws = 0.24676 cjsws = {9.960545E-11*sw_func_psd_nw_cj} cjswgs = {1.47314E-10*sw_func_psd_nw_cj}
+ mjswgs = 0.81 pbs = 0.6587 pbsws = 1
+ pbswgs = 3 xrcrg1 = 12 xrcrg2 = 1
+ rbpb = 50 rbpd = 50 rbps = 50
+ rbdb = 50 rbsb = 50 gbmin = 1E-12
+ tnom = 30 ute = -1.096048 lute = -5.80321E-7
+ wute = -1.734584E-6 pute = 3.311754E-12 kt1 = -0.486836
+ lkt1 = -1.492351E-7 wkt1 = -1.329729E-7 pkt1 = 2.538785E-13
+ kt1l = 0 kt2 = -0.019032 ua1 = 7.780582E-10
+ lua1 = -4.308379E-16 wua1 = -1.574067E-15 pua1 = 3.005287E-21
+ ub1 = -3.361192E-18 lub1 = -5.756547E-25 wub1 = -2.558541E-24
+ pub1 = 4.884894E-30 uc1 = -1.092E-10 at = 2.575737E5
+ lat = -0.203858 wat = 2.13706E-2 pat = -4.08019E-8
+ prt = 0 njs = 1.3632 xtis = 10
+ tpb = 1.671E-3 tpbsw = 0 tpbswg = 0
+ tcj = 9.6E-4 tcjsw = 3E-5 tcjswg = 0
+ tvoff = 0 tvfbsdoff = 0 saref = 3E-6
+ sbref = 3E-6 wlod = 0 ku0 = 7E-8
+ kvsat = 0.4 kvth0 = 3.5E-8 tku0 = 0
+ llodku0 = 0 wlodku0 = 1 llodvth = 0
+ wlodvth = 1 lku0 = 0 wku0 = 0
+ pku0 = 0 lkvth0 = 0 wkvth0 = 6.5E-7
+ pkvth0 = 0 stk2 = 0 lodk2 = 1
+ steta0 = 0 lodeta0 = 1

.model phv_model.19 pmos
+ level = 54 lmin = 8E-7 lmax = 1E-6 wmin = 7E-6
+ wmax = 1.5E-5 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 1.175E-8
+ toxm = 1.175E-8 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 1E23 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {1.2277E-8+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {4.5375E-8-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = -4.7338E-9 dwb = 0 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = -1.124485 lvth0 = 1.074203E-7
+ wvth0 = 8.211076E-7 pvth0 = -5.823705E-13 k1 = 0.590242
+ lk1 = -9.866749E-9 k2 = 2.42311E-2 lk2 = 8.574759E-9
+ wk2 = -2.053956E-8 pk2 = 1.456768E-14 k3 = -2.2405
+ k3b = -0.172 w0 = 0 lpe0 = 0
+ lpeb = 0 vbm = -3 dvtp0 = 0
+ dvtp1 = 0 dvt0 = 4.657 dvt1 = 0.34864
+ dvt2 = -0.030206 dvt0w = -2.2 dvt1w = 1.0163E6
+ dvt2w = 0 vfbsdoff = 0 u0 = 2.16688E-2
+ lu0 = -1.770574E-9 wu0 = -5.028631E-8 pu0 = 3.566556E-14
+ ua = -8.213381E-10 lua = 2.247699E-15 wua = -4.03557E-17
+ pua = 2.862228E-23 ub = 4.622549E-18 lub = -3.399087E-24
+ wub = -6.142872E-24 pub = 4.356832E-30 uc = 6.082696E-12
+ luc = -6.063021E-18 ud = 0 up = 0
+ lp = 1 eu = 1.67 vsat = 8.367108E3
+ lvsat = 3.59353E-2 a0 = 0.824378 la0 = 1.356934E-8
+ wa0 = -4.650489E-7 pa0 = 3.298359E-13 ags = 0.841386
+ lags = -8.529883E-8 wags = -6.925275E-7 pags = 4.911752E-13
+ b0 = 0 b1 = 0 keta = -0.15376
+ lketa = 6.28183E-8 a1 = 0 a2 = 0.5
+ rdsw = 788.47 rdswmin = 0 rdw = 0
+ rdwmin = 0 rsw = 0 rswmin = 0
+ prwb = 0.053538 prwg = 0 wr = 1
+ voff = -9.52546E-2 lvoff = 1.591078E-8 voffl = 0
+ minv = 0 nfactor = 1.014614 lnfactor = 4.665207E-7
+ wnfactor = 4.554915E-6 pnfactor = -3.230573E-12 eta0 = -1.039032E-5
+ leta0 = 4.77441E-11 etab = 7.545356E-4 letab = -6.860615E-10
+ dsub = 1.499307 ldsub = -8.684674E-7 cit = -1.273125E-5
+ lcit = 1.612214E-11 cdsc = 0 cdscb = 0
+ cdscd = 0 pclm = 2.021852 lpclm = -7.444606E-7
+ wpclm = 7.420362E-10 ppclm = -5.262892E-16 pdiblc1 = 0.195862
+ lpdiblc1 = 1.851818E-7 pdiblc2 = -3.36185E-2 lpdiblc2 = 3.193712E-8
+ pdiblcb = -0.025 drout = 0.335842 ldrout = 6.805458E-8
+ pscbe1 = -5.698769E7 lpscbe1 = 324.118516 pscbe2 = 1.828151E-8
+ lpscbe2 = -3.388725E-15 pvag = 0 delta = 0.01
+ fprout = 0 pdits = 0 pditsl = 0
+ pditsd = 0 lambda = 0 vtl = 0
+ lc = 5E-9 xn = 3 alpha0 = 2.471576E-4
+ lalpha0 = -1.63069E-10 alpha1 = 0 beta0 = 67.196894
+ lbeta0 = -1.549723E-5 aigbacc = 0.43 bigbacc = 0.054
+ cigbacc = 0.075 nigbacc = 1 aigbinv = 0.35
+ bigbinv = 0.03 cigbinv = 6E-3 eigbinv = 1.1
+ nigbinv = 3 aigc = 0.43 bigc = 0.054
+ cigc = 0.075 aigsd = 0.43 bigsd = 0.054
+ cigsd = 0.075 dlcig = 0 nigc = 1
+ poxedge = 1 pigcd = 1 ntox = 1
+ toxref = 1.175E-8 agidl = -2.340579E-9 lagidl = 9.717136E-15
+ bgidl = 1.269024E9 lbgidl = 381.772253 cgidl = -171.03
+ lcgidl = 4.90113E-4 egidl = 1.835557 legidl = -9.606931E-7
+ noia = 3E40 noib = 8.53E24 noic = 8.4E7
+ em = 4.1E7 af = 1 ef = 0.88
+ kf = 0 lintnoi = 0 tnoia = 1.5
+ tnoib = 3.5 ntnoi = 1 rnoia = 0.577
+ rnoib = 0.37 xpart = 0 cgso = {1.94171E-10/sw_func_tox_hv_ratio}
+ cgdo = {1.94171E-10/sw_func_tox_hv_ratio} cgbo = {0/sw_func_tox_hv_ratio} ckappas = 0.6
+ cf = 1.2E-11 clc = 1E-7 cle = 0.6
+ dlc = 4.4983E-8 dwc = 0 vfbcv = -0.144689
+ noff = 4 voffcv = 0 acde = 0.401
+ moin = 15.773 cgsl = {9.82591E-12/sw_func_tox_hv_ratio} cgdl = {9.82591E-12/sw_func_tox_hv_ratio}
+ ijthsrev = 0.1 ijthsfwd = 0.1 xjbvs = 1
+ bvs = 12.69 jss = 2.1483E-5 jsws = 4.02E-12
+ cjs = {sw_psd_nw_cj} mjs = 0.33956 mjsws = 0.24676
+ cjsws = {9.960545E-11*sw_func_psd_nw_cj} cjswgs = {1.47314E-10*sw_func_psd_nw_cj} mjswgs = 0.81
+ pbs = 0.6587 pbsws = 1 pbswgs = 3
+ xrcrg1 = 12 xrcrg2 = 1 rbpb = 50
+ rbpd = 50 rbps = 50 rbdb = 50
+ rbsb = 50 gbmin = 1E-12 tnom = 30
+ ute = -2.636771 lute = 8.205817E-7 wute = 8.672919E-6
+ pute = -6.151268E-12 kt1 = -0.677441 lkt1 = 2.407237E-8
+ wkt1 = 6.648644E-7 pkt1 = -4.715551E-13 kt1l = 0
+ kt2 = -0.019032 ua1 = -5.75891E-10 lua1 = 8.002404E-16
+ wua1 = 7.870333E-15 pua1 = -5.582033E-21 ub1 = -5.424862E-18
+ lub1 = 1.300738E-24 wub1 = 1.27927E-23 pub1 = -9.073225E-30
+ uc1 = -1.092E-10 at = 6.304973E4 lat = -2.69868E-2
+ wat = -0.106853 pat = 7.578564E-8 prt = 0
+ njs = 1.3632 xtis = 10 tpb = 1.671E-3
+ tpbsw = 0 tpbswg = 0 tcj = 9.6E-4
+ tcjsw = 3E-5 tcjswg = 0 tvoff = 0
+ tvfbsdoff = 0 saref = 2.81E-6 sbref = 2.81E-6
+ wlod = 0 ku0 = 7E-8 kvsat = 0.4
+ kvth0 = 3.5E-8 tku0 = 0 llodku0 = 0
+ wlodku0 = 1 llodvth = 0 wlodvth = 1
+ lku0 = 0 wku0 = 0 pku0 = 0
+ lkvth0 = 0 wkvth0 = 6.5E-7 pkvth0 = 0
+ stk2 = 0 lodk2 = 1 steta0 = 0
+ lodeta0 = 1

.model phv_model.20 pmos
+ level = 54 lmin = 6E-7 lmax = 8E-7 wmin = 7E-6
+ wmax = 1.5E-5 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 1.175E-8
+ toxm = 1.175E-8 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 1E23 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {1.2277E-8+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {4.5375E-8-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = -4.7338E-9 dwb = 0 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = -0.973029 k1 = 0.57633
+ k2 = 0.036321 k3 = -2.2405 k3b = -0.172
+ w0 = 0 lpe0 = 0 lpeb = 0
+ vbm = -3 dvtp0 = 0 dvtp1 = 0
+ dvt0 = 4.657 dvt1 = 0.34864 dvt2 = -0.030206
+ dvt0w = -2.2 dvt1w = 1.0163E6 dvt2w = 0
+ vfbsdoff = 0 u0 = 1.91724E-2 ua = 2.347784E-9
+ ub = -1.6996E-19 uc = -2.4658E-12 ud = 0
+ up = 0 lp = 1 eu = 1.67
+ vsat = 5.90337E4 a0 = 0.84351 ags = 0.72112
+ b0 = 0 b1 = 0 keta = -0.06519
+ a1 = 0 a2 = 0.5 rdsw = 788.47
+ rdswmin = 0 rdw = 0 rdwmin = 0
+ rsw = 0 rswmin = 0 prwb = 0.053538
+ prwg = 0 wr = 1 voff = -7.28213E-2
+ voffl = 0 minv = 0 nfactor = 1.67238
+ eta0 = 5.6926E-5 etab = -2.1277E-4 dsub = 0.27482
+ cit = 1E-5 cdsc = 0 cdscb = 0
+ cdscd = 0 pclm = 0.972208 pdiblc1 = 0.456957
+ pdiblc2 = 1.14109E-2 pdiblcb = -0.025 drout = 0.431795
+ pscbe1 = 4E8 pscbe2 = 1.350362E-8 pvag = 0
+ delta = 0.01 fprout = 0 pdits = 0
+ pditsl = 0 pditsd = 0 lambda = 0
+ vtl = 0 lc = 5E-9 xn = 3
+ alpha0 = 1.724017E-5 alpha1 = 0 beta0 = 45.34673
+ aigbacc = 0.43 bigbacc = 0.054 cigbacc = 0.075
+ nigbacc = 1 aigbinv = 0.35 bigbinv = 0.03
+ cigbinv = 6E-3 eigbinv = 1.1 nigbinv = 3
+ aigc = 0.43 bigc = 0.054 cigc = 0.075
+ aigsd = 0.43 bigsd = 0.054 cigsd = 0.075
+ dlcig = 0 nigc = 1 poxedge = 1
+ pigcd = 1 ntox = 1 toxref = 1.175E-8
+ agidl = 1.136E-8 bgidl = 1.8073E9 cgidl = 520
+ egidl = 0.481037 noia = 3E40 noib = 8.53E24
+ noic = 8.4E7 em = 4.1E7 af = 1
+ ef = 0.88 kf = 0 lintnoi = 0
+ tnoia = 1.5 tnoib = 3.5 ntnoi = 1
+ rnoia = 0.577 rnoib = 0.37 xpart = 0
+ cgso = {1.94171E-10/sw_func_tox_hv_ratio} cgdo = {1.94171E-10/sw_func_tox_hv_ratio} cgbo = {0/sw_func_tox_hv_ratio}
+ ckappas = 0.6 cf = 1.2E-11 clc = 1E-7
+ cle = 0.6 dlc = 4.4983E-8 dwc = 0
+ vfbcv = -0.144689 noff = 4 voffcv = 0
+ acde = 0.401 moin = 15.773 cgsl = {9.82591E-12/sw_func_tox_hv_ratio}
+ cgdl = {9.82591E-12/sw_func_tox_hv_ratio} ijthsrev = 0.1 ijthsfwd = 0.1
+ xjbvs = 1 bvs = 12.69 jss = 2.1483E-5
+ jsws = 4.02E-12 cjs = {sw_psd_nw_cj} mjs = 0.33956
+ mjsws = 0.24676 cjsws = {9.960545E-11*sw_func_psd_nw_cj} cjswgs = {1.47314E-10*sw_func_psd_nw_cj}
+ mjswgs = 0.81 pbs = 0.6587 pbsws = 1
+ pbswgs = 3 xrcrg1 = 12 xrcrg2 = 1
+ rbpb = 50 rbpd = 50 rbps = 50
+ rbdb = 50 rbsb = 50 gbmin = 1E-12
+ tnom = 30 ute = -1.4798 kt1 = -0.6435
+ kt1l = 0 kt2 = -0.019032 ua1 = 5.524E-10
+ ub1 = -3.5909E-18 uc1 = -1.092E-10 at = 2.5E4
+ prt = 0 njs = 1.3632 xtis = 10
+ tpb = 1.671E-3 tpbsw = 0 tpbswg = 0
+ tcj = 9.6E-4 tcjsw = 3E-5 tcjswg = 0
+ tvoff = 0 tvfbsdoff = 0 saref = 2.41E-6
+ sbref = 2.41E-6 wlod = 0 ku0 = 7E-8
+ kvsat = 0.4 kvth0 = 3.5E-8 tku0 = 0
+ llodku0 = 0 wlodku0 = 1 llodvth = 0
+ wlodvth = 1 lku0 = 0 wku0 = 0
+ pku0 = 0 lkvth0 = 0 wkvth0 = 6.5E-7
+ pkvth0 = 0 stk2 = 0 lodk2 = 1
+ steta0 = 0 lodeta0 = 1

.model phv_model.21 pmos
+ level = 54 lmin = 5E-7 lmax = 6E-7 wmin = 7E-6
+ wmax = 1.5E-5 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 1.175E-8
+ toxm = 1.175E-8 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 1E23 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {1.2277E-8+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {4.5375E-8-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = -4.7338E-9 dwb = 0 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = -0.753132 lvth0 = -1.119827E-7
+ wvth0 = -6.697923E-7 pvth0 = 3.410917E-13 k1 = 0.487482
+ lk1 = 4.524593E-8 k2 = 3.09905E-2 lk2 = 2.71455E-9
+ wk2 = -3.48416E-8 pk2 = 1.774308E-14 k3 = -2.2405
+ k3b = -0.172 w0 = 0 lpe0 = 0
+ lpeb = 0 vbm = -3 dvtp0 = 0
+ dvtp1 = 0 dvt0 = 4.657 dvt1 = 0.34864
+ dvt2 = -0.030206 dvt0w = -2.2 dvt1w = 1.0163E6
+ dvt2w = 0 vfbsdoff = 0 u0 = 1.10187E-2
+ lu0 = 4.152256E-9 wu0 = 4.558798E-8 pu0 = -2.321568E-14
+ ua = 3.12154E-9 lua = -3.940357E-16 wua = -4.216314E-17
+ pua = 2.147158E-23 ub = -3.876447E-18 lub = 1.887528E-24
+ wub = 9.047059E-24 pub = -4.607215E-30 uc = 9.057452E-12
+ luc = -5.868216E-18 ud = 0 up = 0
+ lp = 1 eu = 1.67 vsat = 3.932107E4
+ lvsat = 1.00387E-2 wvsat = 2.57571E-2 pvsat = -1.311682E-8
+ a0 = 0.368248 la0 = 2.420272E-7 ags = -1.443321
+ lags = 1.102242E-6 b0 = 0 b1 = 0
+ keta = 1.94429E-2 lketa = -4.30993E-8 a1 = 0
+ a2 = 0.5 rdsw = 788.47 rdswmin = 0
+ rdw = 0 rdwmin = 0 rsw = 0
+ rswmin = 0 prwb = 0.053538 prwg = 0
+ wr = 1 voff = 4.46966E-2 lvoff = -5.984601E-8
+ voffl = 0 minv = 0 nfactor = 1.816498
+ lnfactor = -7.339218E-8 wnfactor = -3.957621E-6 pnfactor = 2.015418E-12
+ eta0 = -0.241472 leta0 = 1.229986E-7 weta0 = -5.989335E-7
+ peta0 = 3.050069E-13 etab = 1.46738E-2 letab = -7.580997E-9
+ dsub = 0.254971 ldsub = 1.010791E-8 cit = 3.04625E-5
+ lcit = -1.042053E-11 cdsc = 0 cdscb = 0
+ cdscd = 0 pclm = -0.518953 lpclm = 7.593738E-7
+ wpclm = -1.715361E-9 ppclm = 8.735475E-16 pdiblc1 = 1.123736
+ lpdiblc1 = -3.39557E-7 pdiblc2 = 3.84625E-2 lpdiblc2 = -1.377603E-8
+ pdiblcb = -0.025 drout = -1.482714 ldrout = 9.749638E-7
+ pscbe1 = 5.52896E8 lpscbe1 = -77.86227 pscbe2 = 9.480217E-9
+ lpscbe2 = 2.048916E-15 pvag = 0 delta = 0.01
+ fprout = 0 pdits = 0 pditsl = 0
+ pditsd = 0 lambda = 0 vtl = 0
+ lc = 5E-9 xn = 3 alpha0 = -3.097308E-4
+ lalpha0 = 1.6651E-10 alpha1 = 0 beta0 = 7.131861
+ lbeta0 = 1.946092E-5 aigbacc = 0.43 bigbacc = 0.054
+ cigbacc = 0.075 nigbacc = 1 aigbinv = 0.35
+ bigbinv = 0.03 cigbinv = 6E-3 eigbinv = 1.1
+ nigbinv = 3 aigc = 0.43 bigc = 0.054
+ cigc = 0.075 aigsd = 0.43 bigsd = 0.054
+ cigsd = 0.075 dlcig = 0 nigc = 1
+ poxedge = 1 pigcd = 1 ntox = 1
+ toxref = 1.175E-8 agidl = -1.046062E-8 lagidl = 1.111215E-14
+ wagidl = 1.853231E-13 pagidl = -9.437578E-20 bgidl = 2.353562E9
+ lbgidl = -278.183739 wbgidl = 3.329189E3 pbgidl = -1.69539E-3
+ cgidl = 842.951128 lcgidl = -1.644629E-4 wcgidl = 7.624538E-3
+ pcgidl = -3.882796E-9 egidl = -0.272932 legidl = 3.839585E-7
+ noia = 3E40 noib = 8.53E24 noic = 8.4E7
+ em = 4.1E7 af = 1 ef = 0.88
+ kf = 0 lintnoi = 0 tnoia = 1.5
+ tnoib = 3.5 ntnoi = 1 rnoia = 0.577
+ rnoib = 0.37 xpart = 0 cgso = {1.94171E-10/sw_func_tox_hv_ratio}
+ cgdo = {1.94171E-10/sw_func_tox_hv_ratio} cgbo = {0/sw_func_tox_hv_ratio} ckappas = 0.6
+ cf = 1.2E-11 clc = 1E-7 cle = 0.6
+ dlc = 4.4983E-8 dwc = 0 vfbcv = -0.144689
+ noff = 4 voffcv = 0 acde = 0.401
+ moin = 15.773 cgsl = {9.82591E-12/sw_func_tox_hv_ratio} cgdl = {9.82591E-12/sw_func_tox_hv_ratio}
+ ijthsrev = 0.1 ijthsfwd = 0.1 xjbvs = 1
+ bvs = 12.69 jss = 2.1483E-5 jsws = 4.02E-12
+ cjs = {sw_psd_nw_cj} mjs = 0.33956 mjsws = 0.24676
+ cjsws = {9.960545E-11*sw_func_psd_nw_cj} cjswgs = {1.47314E-10*sw_func_psd_nw_cj} mjswgs = 0.81
+ pbs = 0.6587 pbsws = 1 pbswgs = 3
+ xrcrg1 = 12 xrcrg2 = 1 rbpb = 50
+ rbpd = 50 rbps = 50 rbdb = 50
+ rbsb = 50 gbmin = 1E-12 tnom = 30
+ ute = -1.919334 lute = 2.238329E-7 kt1 = -0.807282
+ lkt1 = 8.340591E-8 kt1l = 0 kt2 = -0.019032
+ ua1 = 5.524E-10 ub1 = -9.446858E-18 lub1 = 2.982147E-24
+ uc1 = -3.862786E-10 luc1 = 1.411023E-16 at = 5.36475E4
+ lat = -1.45887E-2 prt = 0 njs = 1.3632
+ xtis = 10 tpb = 1.671E-3 tpbsw = 0
+ tpbswg = 0 tcj = 9.6E-4 tcjsw = 3E-5
+ tcjswg = 0 tvoff = 0 tvfbsdoff = 0
+ saref = 2.41E-6 sbref = 2.41E-6 wlod = 0
+ ku0 = 7E-8 kvsat = 0.4 kvth0 = 3.5E-8
+ tku0 = 0 llodku0 = 0 wlodku0 = 1
+ llodvth = 0 wlodvth = 1 lku0 = 0
+ wku0 = 0 pku0 = 0 lkvth0 = 0
+ wkvth0 = 6.5E-7 pkvth0 = 0 stk2 = 0
+ lodk2 = 1 steta0 = 0 lodeta0 = 1

.model phv_model.22 pmos
+ level = 54 lmin = 8E-6 lmax = 2.02E-5 wmin = 3E-6
+ wmax = 7E-6 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 1.175E-8
+ toxm = 1.175E-8 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 1E23 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {1.2277E-8+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {4.5375E-8-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = -4.7338E-9 dwb = 0 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = -1.029992 wvth0 = 1.322829E-7
+ k1 = 0.59521 k2 = 2.55231E-2 wk2 = -1.693094E-9
+ k3 = -2.2405 k3b = -0.172 w0 = 0
+ lpe0 = 0 lpeb = 0 vbm = -3
+ dvtp0 = 0 dvtp1 = 0 dvt0 = 4.657
+ dvt1 = 0.34864 dvt2 = -0.030206 dvt0w = -2.2
+ dvt1w = 1.0163E6 dvt2w = 0 vfbsdoff = 0
+ u0 = 2.18988E-2 wu0 = -6.369729E-9 ua = 2.746957E-9
+ wua = -2.967748E-16 ub = -1.576849E-19 wub = -1.224549E-25
+ uc = -3.9972E-11 ud = 0 up = 0
+ lp = 1 eu = 1.67 vsat = 2E5
+ a0 = 0.716278 wa0 = 1.258797E-6 ags = 0.115609
+ wags = 1.301892E-7 b0 = 0 b1 = 0
+ keta = -7.9259E-3 a1 = 0 a2 = 0.5
+ rdsw = 788.47 rdswmin = 0 rdw = 0
+ rdwmin = 0 rsw = 0 rswmin = 0
+ prwb = 0.053538 prwg = 0 wr = 1
+ voff = -9.32047E-2 voffl = 0 minv = 0
+ nfactor = 1.73965 eta0 = 0.08 etab = -0.07
+ dsub = 0.56 cit = 1E-5 cdsc = 0
+ cdscb = 0 cdscd = 0 pclm = 8.35312E-2
+ pdiblc1 = 0.39 pdiblc2 = 2.940788E-3 pdiblcb = -0.025
+ drout = 0.56 pscbe1 = 3.337128E8 pscbe2 = 1.500096E-8
+ pvag = 0 delta = 0.01 fprout = 0
+ pdits = 0 pditsl = 0 pditsd = 0
+ lambda = 0 vtl = 0 lc = 5E-9
+ xn = 3 alpha0 = 5.066719E-5 alpha1 = 0
+ beta0 = 38.266046 aigbacc = 0.43 bigbacc = 0.054
+ cigbacc = 0.075 nigbacc = 1 aigbinv = 0.35
+ bigbinv = 0.03 cigbinv = 6E-3 eigbinv = 1.1
+ nigbinv = 3 aigc = 0.43 bigc = 0.054
+ cigc = 0.075 aigsd = 0.43 bigsd = 0.054
+ cigsd = 0.075 dlcig = 0 nigc = 1
+ poxedge = 1 pigcd = 1 ntox = 1
+ toxref = 1.175E-8 agidl = 1.854207E-9 wagidl = 3.844512E-14
+ bgidl = 1.651886E9 wbgidl = 368.402366 cgidl = 476.84155
+ wcgidl = 1.55663E-3 egidl = 0.693508 noia = 3E40
+ noib = 8.53E24 noic = 8.4E7 em = 4.1E7
+ af = 1 ef = 0.88 kf = 0
+ lintnoi = 0 tnoia = 1.5 tnoib = 3.5
+ ntnoi = 1 rnoia = 0.577 rnoib = 0.37
+ xpart = 0 cgso = {1.94171E-10/sw_func_tox_hv_ratio} cgdo = {1.94171E-10/sw_func_tox_hv_ratio}
+ cgbo = {0/sw_func_tox_hv_ratio} ckappas = 0.6 cf = 1.2E-11
+ clc = 1E-7 cle = 0.6 dlc = 4.4983E-8
+ dwc = 0 vfbcv = -0.144689 noff = 4
+ voffcv = 0 acde = 0.401 moin = 15.773
+ cgsl = {9.82591E-12/sw_func_tox_hv_ratio} cgdl = {9.82591E-12/sw_func_tox_hv_ratio} ijthsrev = 0.1
+ ijthsfwd = 0.1 xjbvs = 1 bvs = 12.69
+ jss = 2.1483E-5 jsws = 4.02E-12 cjs = {sw_psd_nw_cj}
+ mjs = 0.33956 mjsws = 0.24676 cjsws = {9.960545E-11*sw_func_psd_nw_cj}
+ cjswgs = {1.47314E-10*sw_func_psd_nw_cj} mjswgs = 0.81 pbs = 0.6587
+ pbsws = 1 pbswgs = 3 xrcrg1 = 12
+ xrcrg2 = 1 rbpb = 50 rbpd = 50
+ rbps = 50 rbdb = 50 rbsb = 50
+ gbmin = 1E-12 tnom = 30 ute = -1.275044
+ wute = -7.767582E-7 kt1 = -0.576 kt1l = 0
+ kt2 = -0.019032 ua1 = 1.215706E-9 wua1 = -3.551523E-15
+ ub1 = -2.759903E-18 wub1 = -2.686224E-24 uc1 = -1.092E-10
+ at = 4.160154E5 wat = 9.75488E-2 prt = 0
+ njs = 1.3632 xtis = 10 tpb = 1.671E-3
+ tpbsw = 0 tpbswg = 0 tcj = 9.6E-4
+ tcjsw = 3E-5 tcjswg = 0 tvoff = 0
+ tvfbsdoff = 0 saref = 3E-6 sbref = 3E-6
+ wlod = 0 ku0 = 7E-8 kvsat = 0.4
+ kvth0 = 3.5E-8 tku0 = 0 llodku0 = 0
+ wlodku0 = 1 llodvth = 0 wlodvth = 1
+ lku0 = 0 wku0 = 0 pku0 = 0
+ lkvth0 = 0 wkvth0 = 6.5E-7 pkvth0 = 0
+ stk2 = 0 lodk2 = 1 steta0 = 0
+ lodeta0 = 1

.model phv_model.23 pmos
+ level = 54 lmin = 4E-6 lmax = 8E-6 wmin = 3E-6
+ wmax = 7E-6 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 1.175E-8
+ toxm = 1.175E-8 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 1E23 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {1.2277E-8+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {4.5375E-8-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = -4.7338E-9 dwb = 0 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = -1.037268 lvth0 = 5.754762E-8
+ wvth0 = 1.46496E-7 pvth0 = -1.124152E-13 k1 = 0.604152
+ lk1 = -7.072775E-8 k2 = 2.30493E-2 lk2 = 1.956599E-8
+ wk2 = 1.745075E-9 pk2 = -2.719334E-14 k3 = -2.2405
+ k3b = -0.172 w0 = 0 lpe0 = 0
+ lpeb = 0 vbm = -3 dvtp0 = 0
+ dvtp1 = 0 dvt0 = 4.657 dvt1 = 0.34864
+ dvt2 = -0.030206 dvt0w = -2.2 dvt1w = 1.0163E6
+ dvt2w = 0 vfbsdoff = 0 u0 = 2.12187E-2
+ lu0 = 5.379018E-9 wu0 = -6.745493E-9 pu0 = 2.972015E-15
+ ua = 2.533417E-9 lua = 1.688945E-15 wua = -5.835026E-16
+ pua = 2.267801E-21 ub = 3.522753E-20 lub = -1.525792E-24
+ wub = 3.717185E-25 pub = -3.908541E-30 uc = -5.157563E-11
+ luc = 9.177602E-17 ud = 0 up = 0
+ lp = 1 eu = 1.67 vsat = 3.158234E5
+ lvsat = -0.916076 wvsat = -0.126269 pvsat = 9.986934E-7
+ a0 = 0.560839 la0 = 1.229406E-6 wa0 = 2.481182E-6
+ pa0 = -9.668146E-12 ags = 0.066077 lags = 3.917645E-7
+ wags = 3.046991E-7 pags = -1.380242E-12 b0 = 0
+ b1 = 0 keta = -4.956727E-3 lketa = -2.348393E-8
+ a1 = 0 a2 = 0.5 rdsw = 788.47
+ rdswmin = 0 rdw = 0 rdwmin = 0
+ rsw = 0 rswmin = 0 prwb = 0.053538
+ prwg = 0 wr = 1 voff = -9.47765E-2
+ lvoff = 1.243193E-8 voffl = 0 minv = 0
+ nfactor = 1.771232 lnfactor = -2.437187E-7 wnfactor = -1.119698E-7
+ pnfactor = 8.675397E-13 eta0 = 0.08 etab = -0.07
+ dsub = 0.56 cit = 1E-5 cdsc = 0
+ cdscb = 0 cdscd = 0 pclm = -0.648319
+ lpclm = 5.788389E-6 pdiblc1 = 0.39 pdiblc2 = 4.554123E-3
+ lpdiblc2 = -1.276027E-8 pdiblcb = -0.025 drout = 0.56
+ pscbe1 = 5.621233E8 lpscbe1 = -1.806556E3 pscbe2 = -1.531739E-8
+ lpscbe2 = 2.397954E-13 pvag = 0 delta = 0.01
+ fprout = 0 pdits = 0 pditsl = 0
+ pditsd = 0 lambda = 0 vtl = 0
+ lc = 5E-9 xn = 3 alpha0 = 7.815322E-5
+ lalpha0 = -2.173939E-10 alpha1 = 0 beta0 = 39.140288
+ lbeta0 = -6.9146E-6 aigbacc = 0.43 bigbacc = 0.054
+ cigbacc = 0.075 nigbacc = 1 aigbinv = 0.35
+ bigbinv = 0.03 cigbinv = 6E-3 eigbinv = 1.1
+ nigbinv = 3 aigc = 0.43 bigc = 0.054
+ cigc = 0.075 aigsd = 0.43 bigsd = 0.054
+ cigsd = 0.075 dlcig = 0 nigc = 1
+ poxedge = 1 pigcd = 1 ntox = 1
+ toxref = 1.175E-8 agidl = -3.495344E-9 lagidl = 4.231094E-14
+ wagidl = 6.99926E-14 pagidl = -2.495169E-19 bgidl = 1.319764E9
+ lbgidl = 2.626835E3 wbgidl = 1.10624E3 pbgidl = -5.835738E-3
+ cgidl = 635.28944 lcgidl = -1.253204E-3 wcgidl = 2.073876E-3
+ pcgidl = -4.091033E-9 egidl = 1.209319 legidl = -4.079675E-6
+ noia = 3E40 noib = 8.53E24 noic = 8.4E7
+ em = 4.1E7 af = 1 ef = 0.88
+ kf = 0 lintnoi = 0 tnoia = 1.5
+ tnoib = 3.5 ntnoi = 1 rnoia = 0.577
+ rnoib = 0.37 xpart = 0 cgso = {1.94171E-10/sw_func_tox_hv_ratio}
+ cgdo = {1.94171E-10/sw_func_tox_hv_ratio} cgbo = {0/sw_func_tox_hv_ratio} ckappas = 0.6
+ cf = 1.2E-11 clc = 1E-7 cle = 0.6
+ dlc = 4.4983E-8 dwc = 0 vfbcv = -0.144689
+ noff = 4 voffcv = 0 acde = 0.401
+ moin = 15.773 cgsl = {9.82591E-12/sw_func_tox_hv_ratio} cgdl = {9.82591E-12/sw_func_tox_hv_ratio}
+ ijthsrev = 0.1 ijthsfwd = 0.1 xjbvs = 1
+ bvs = 12.69 jss = 2.1483E-5 jsws = 4.02E-12
+ cjs = {sw_psd_nw_cj} mjs = 0.33956 mjsws = 0.24676
+ cjsws = {9.960545E-11*sw_func_psd_nw_cj} cjswgs = {1.47314E-10*sw_func_psd_nw_cj} mjswgs = 0.81
+ pbs = 0.6587 pbsws = 1 pbswgs = 3
+ xrcrg1 = 12 xrcrg2 = 1 rbpb = 50
+ rbpd = 50 rbps = 50 rbdb = 50
+ rbsb = 50 gbmin = 1E-12 tnom = 30
+ ute = -1.000364 lute = -2.17251E-6 wute = -1.535894E-6
+ pute = 6.004193E-12 kt1 = -0.592112 lkt1 = 1.311576E-7
+ wkt1 = 4.794031E-8 pkt1 = -3.902525E-13 kt1l = 0
+ kt2 = -0.019032 ua1 = 2.382237E-9 lua1 = -9.22638E-15
+ wua1 = -7.022472E-15 pua1 = 2.74526E-20 ub1 = -1.893735E-18
+ lub1 = -6.850738E-24 wub1 = -4.999128E-24 pub1 = 1.829334E-29
+ uc1 = -1.092E-10 at = 6.805457E5 lat = -2.092236
+ wat = -5.23006E-2 pat = 1.185196E-6 prt = 0
+ njs = 1.3632 xtis = 10 tpb = 1.671E-3
+ tpbsw = 0 tpbswg = 0 tcj = 9.6E-4
+ tcjsw = 3E-5 tcjswg = 0 tvoff = 0
+ tvfbsdoff = 0 saref = 3E-6 sbref = 3E-6
+ wlod = 0 ku0 = 7E-8 kvsat = 0.4
+ kvth0 = 3.5E-8 tku0 = 0 llodku0 = 0
+ wlodku0 = 1 llodvth = 0 wlodvth = 1
+ lku0 = 0 wku0 = 0 pku0 = 0
+ lkvth0 = 0 wkvth0 = 6.5E-7 pkvth0 = 0
+ stk2 = 0 lodk2 = 1 steta0 = 0
+ lodeta0 = 1

.model phv_model.24 pmos
+ level = 54 lmin = 2E-6 lmax = 4E-6 wmin = 3E-6
+ wmax = 7E-6 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 1.175E-8
+ toxm = 1.175E-8 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 1E23 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {1.2277E-8+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {4.5375E-8-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = -4.7338E-9 dwb = 0 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = -1.005773 lvth0 = -6.557502E-8
+ wvth0 = 1.020938E-7 pvth0 = 6.11644E-14 k1 = 0.602594
+ lk1 = -6.463595E-8 k2 = 2.79207E-2 lk2 = 5.224713E-10
+ wk2 = -7.593627E-9 pk2 = 9.313982E-15 k3 = -2.2405
+ k3b = -0.172 w0 = 0 lpe0 = 0
+ lpeb = 0 vbm = -3 dvtp0 = 0
+ dvtp1 = 0 dvt0 = 4.657 dvt1 = 0.34864
+ dvt2 = -0.030206 dvt0w = -2.2 dvt1w = 1.0163E6
+ dvt2w = 0 vfbsdoff = 0 u0 = 2.17997E-2
+ lu0 = 3.107763E-9 wu0 = -6.008126E-9 pu0 = 8.94607E-17
+ ua = 3.313609E-9 lua = -1.361023E-15 wua = 1.791108E-18
+ pua = -2.025801E-23 ub = -1.317733E-18 lub = 3.76327E-24
+ wub = -9.923132E-25 pub = 1.4238E-30 uc = -5.492301E-11
+ luc = 1.048618E-16 ud = 0 up = 0
+ lp = 1 eu = 1.67 vsat = 6.254339E4
+ lvsat = 7.40586E-2 wvsat = 0.153472 pvsat = -9.488256E-8
+ a0 = 0.820219 la0 = 2.154241E-7 wa0 = 2.443581E-8
+ pa0 = -6.411156E-14 ags = 0.128532 lags = 1.476137E-7
+ wags = -5.039662E-8 pags = 7.915723E-15 b0 = 0
+ b1 = 0 keta = -5.087328E-3 lketa = -2.297338E-8
+ a1 = 0 a2 = 0.5 rdsw = 788.47
+ rdswmin = 0 rdw = 0 rdwmin = 0
+ rsw = 0 rswmin = 0 prwb = 0.053538
+ prwg = 0 wr = 1 voff = -0.064087
+ lvoff = -1.075408E-7 voffl = 0 minv = 0
+ nfactor = 2.048398 lnfactor = -1.32723E-6 wnfactor = 7.510539E-7
+ pnfactor = -2.506236E-12 eta0 = 1.90949E-2 leta0 = 2.380932E-7
+ etab = -0.122401 letab = 2.048497E-7 dsub = 0.814742
+ ldsub = -9.958489E-7 cit = 1E-5 cdsc = 0
+ cdscb = 0 cdscd = 0 pclm = 1.048765
+ lpclm = -8.459384E-7 ppclm = -1.587831E-17 pdiblc1 = 0.581562
+ lpdiblc1 = -7.488642E-7 pdiblc2 = -1.133342E-3 lpdiblc2 = 9.473451E-9
+ pdiblcb = 0.165925 lpdiblcb = -7.463736E-7 drout = 0.139965
+ ldrout = 1.642022E-6 pscbe1 = -1.561704E8 lpscbe1 = 1.001434E3
+ pscbe2 = 7.607469E-8 lpscbe2 = -1.174791E-13 pvag = 0
+ delta = 0.01 fprout = 0 pdits = 0
+ pditsl = 0 pditsd = 0 lambda = 0
+ vtl = 0 lc = 5E-9 xn = 3
+ alpha0 = 4.406319E-5 lalpha0 = -8.412745E-11 alpha1 = -9.54625E-11
+ lalpha1 = 3.731868E-16 beta0 = 70.183411 lbeta0 = -1.282699E-4
+ aigbacc = 0.43 bigbacc = 0.054 cigbacc = 0.075
+ nigbacc = 1 aigbinv = 0.35 bigbinv = 0.03
+ cigbinv = 6E-3 eigbinv = 1.1 nigbinv = 3
+ aigc = 0.43 bigc = 0.054 cigc = 0.075
+ aigsd = 0.43 bigsd = 0.054 cigsd = 0.075
+ dlcig = 0 nigc = 1 poxedge = 1
+ pigcd = 1 ntox = 1 toxref = 1.175E-8
+ agidl = 8.985284E-9 lagidl = -6.478956E-15 wagidl = 1.47796E-15
+ pagidl = 1.832395E-20 bgidl = 2.728323E9 lbgidl = -2.879575E3
+ wbgidl = -755.585795 pbgidl = 1.442602E-3 cgidl = 167.86109
+ lcgidl = 5.740903E-4 wcgidl = 2.008134E-3 pcgidl = -3.83403E-9
+ egidl = -1.585323 legidl = 6.845277E-6 noia = 3E40
+ noib = 8.53E24 noic = 8.4E7 em = 4.1E7
+ af = 1 ef = 0.88 kf = 0
+ lintnoi = 0 tnoia = 1.5 tnoib = 3.5
+ ntnoi = 1 rnoia = 0.577 rnoib = 0.37
+ xpart = 0 cgso = {1.94171E-10/sw_func_tox_hv_ratio} cgdo = {1.94171E-10/sw_func_tox_hv_ratio}
+ cgbo = {0/sw_func_tox_hv_ratio} ckappas = 0.6 cf = 1.2E-11
+ clc = 1E-7 cle = 0.6 dlc = 4.4983E-8
+ dwc = 0 vfbcv = -0.144689 noff = 4
+ voffcv = 0 acde = 0.401 moin = 15.773
+ cgsl = {9.82591E-12/sw_func_tox_hv_ratio} cgdl = {9.82591E-12/sw_func_tox_hv_ratio} ijthsrev = 0.1
+ ijthsfwd = 0.1 xjbvs = 1 bvs = 12.69
+ jss = 2.1483E-5 jsws = 4.02E-12 cjs = {sw_psd_nw_cj}
+ mjs = 0.33956 mjsws = 0.24676 cjsws = {9.960545E-11*sw_func_psd_nw_cj}
+ cjswgs = {1.47314E-10*sw_func_psd_nw_cj} mjswgs = 0.81 pbs = 0.6587
+ pbsws = 1 pbswgs = 3 xrcrg1 = 12
+ xrcrg2 = 1 rbpb = 50 rbpd = 50
+ rbps = 50 rbdb = 50 rbsb = 50
+ gbmin = 1E-12 tnom = 30 ute = -1.74048
+ lute = 7.20789E-7 wute = 2.466756E-7 pute = -9.643166E-13
+ kt1 = -0.559516 lkt1 = 3.731868E-9 wkt1 = -5.188766E-8
+ kt1l = 0 kt2 = -0.019032 ua1 = -4.841455E-10
+ lua1 = 1.979024E-15 ub1 = -3.956417E-18 lub1 = 1.212801E-24
+ wub1 = 1.649319E-24 pub1 = -7.697106E-30 uc1 = -1.092E-10
+ at = 1.549987E5 lat = -3.77416E-2 wat = 0.386697
+ pat = -5.309551E-7 prt = 0 njs = 1.3632
+ xtis = 10 tpb = 1.671E-3 tpbsw = 0
+ tpbswg = 0 tcj = 9.6E-4 tcjsw = 3E-5
+ tcjswg = 0 tvoff = 0 tvfbsdoff = 0
+ saref = 3E-6 sbref = 3E-6 wlod = 0
+ ku0 = 7E-8 kvsat = 0.4 kvth0 = 3.5E-8
+ tku0 = 0 llodku0 = 0 wlodku0 = 1
+ llodvth = 0 wlodvth = 1 lku0 = 0
+ wku0 = 0 pku0 = 0 lkvth0 = 0
+ wkvth0 = 6.5E-7 pkvth0 = 0 stk2 = 0
+ lodk2 = 1 steta0 = 0 lodeta0 = 1

.model phv_model.25 pmos
+ level = 54 lmin = 1E-6 lmax = 2E-6 wmin = 3E-6
+ wmax = 7E-6 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 1.175E-8
+ toxm = 1.175E-8 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 1E23 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {1.2277E-8+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {4.5375E-8-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = -4.7338E-9 dwb = 0 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = -1.078862 lvth0 = 7.397092E-8
+ wvth0 = 1.479011E-7 pvth0 = -2.629325E-14 k1 = 0.559056
+ lk1 = 1.848825E-8 k2 = 2.31678E-2 lk2 = 9.596968E-9
+ wk2 = -6.898081E-10 pk2 = -3.867134E-15 k3 = -2.2405
+ k3b = -0.172 w0 = 0 lpe0 = 0
+ lpeb = 0 vbm = -3 dvtp0 = 0
+ dvtp1 = 0 dvt0 = 4.657 dvt1 = 0.34864
+ dvt2 = -0.030206 dvt0w = -2.2 dvt1w = 1.0163E6
+ dvt2w = 0 vfbsdoff = 0 u0 = 2.75761E-2
+ lu0 = -7.920906E-9 wu0 = -6.758969E-9 pu0 = 1.523009E-15
+ ua = 3.465241E-9 lua = -1.650525E-15 wua = -1.332353E-17
+ pua = 8.59961E-24 ub = 5.787865E-19 lub = 1.423395E-25
+ wub = -1.86427E-25 pub = -1.148382E-31 uc = 5.323295E-13
+ luc = -1.01635E-18 ud = 0 up = 0
+ lp = 1 eu = 1.67 vsat = 1.499265E5
+ lvsat = -9.27776E-2 wvsat = 0.198133 pvsat = -1.801524E-7
+ a0 = 1.046318 la0 = -2.162538E-7 wa0 = -1.199319E-7
+ pa0 = 2.115224E-13 ags = -0.282543 lags = 9.324585E-7
+ wags = 2.1075E-8 pags = -1.285415E-13 b0 = 0
+ b1 = 0 keta = 4.43017E-2 lketa = -1.172693E-7
+ a1 = 0 a2 = 0.5 rdsw = 788.47
+ rdswmin = 0 rdw = 0 rdwmin = 0
+ rsw = 0 rswmin = 0 prwb = 0.053538
+ prwg = 0 wr = 1 voff = -0.1592
+ lvoff = 7.405273E-8 voffl = 0 minv = 0
+ nfactor = 1.066289 lnfactor = 5.478611E-7 wnfactor = -1.088138E-6
+ pnfactor = 1.005242E-12 eta0 = 0.280418 leta0 = -2.608385E-7
+ weta0 = -4.120026E-8 peta0 = 7.866159E-14 etab = -2.88449E-2
+ letab = 2.622727E-8 dsub = -0.100903 ldsub = 7.523465E-7
+ wdsub = 1.156686E-6 pdsub = -2.208403E-12 cit = 1.454625E-5
+ lcit = -8.679928E-12 cdsc = 0 cdscb = 0
+ cdscd = 0 pclm = 6.24863E-2 lpclm = 1.037114E-6
+ ppclm = 7.38625E-18 pdiblc1 = -1.786113E-3 lpdiblc1 = 3.648934E-7
+ pdiblc2 = 5.940119E-3 lpdiblc2 = -4.031554E-9 pdiblcb = -0.40685
+ lpdiblcb = 3.471971E-7 drout = 1.535831 ldrout = -1.023035E-6
+ pscbe1 = 4.309632E8 lpscbe1 = -119.550868 pscbe2 = 1.454314E-8
+ pvag = 0 delta = 0.01 fprout = 0
+ pdits = 0 pditsl = 0 pditsd = 0
+ lambda = 0 vtl = 0 lc = 5E-9
+ xn = 3 alpha0 = -6.165893E-5 lalpha0 = 1.177225E-10
+ alpha1 = 1.90925E-10 lalpha1 = -1.735986E-16 beta0 = -39.873797
+ lbeta0 = 8.18568E-5 aigbacc = 0.43 bigbacc = 0.054
+ cigbacc = 0.075 nigbacc = 1 aigbinv = 0.35
+ bigbinv = 0.03 cigbinv = 6E-3 eigbinv = 1.1
+ nigbinv = 3 aigc = 0.43 bigc = 0.054
+ cigc = 0.075 aigsd = 0.43 bigsd = 0.054
+ cigsd = 0.075 dlcig = 0 nigc = 1
+ poxedge = 1 pigcd = 1 ntox = 1
+ toxref = 1.175E-8 agidl = 1.50997E-9 lagidl = 7.793286E-15
+ wagidl = 3.214785E-14 pagidl = -4.023255E-20 bgidl = 7.092315E8
+ lbgidl = 975.375768 wbgidl = 590.207443 pbgidl = -1.126854E-3
+ cgidl = 933.323638 lcgidl = -8.873691E-4 wcgidl = -2.604273E-3
+ pcgidl = 4.972208E-9 egidl = 3.110213 legidl = -2.119675E-6
+ noia = 3E40 noib = 8.53E24 noic = 8.4E7
+ em = 4.1E7 af = 1 ef = 0.88
+ kf = 0 lintnoi = 0 tnoia = 1.5
+ tnoib = 3.5 ntnoi = 1 rnoia = 0.577
+ rnoib = 0.37 xpart = 0 cgso = {1.94171E-10/sw_func_tox_hv_ratio}
+ cgdo = {1.94171E-10/sw_func_tox_hv_ratio} cgbo = {0/sw_func_tox_hv_ratio} ckappas = 0.6
+ cf = 1.2E-11 clc = 1E-7 cle = 0.6
+ dlc = 4.4983E-8 dwc = 0 vfbcv = -0.144689
+ noff = 4 voffcv = 0 acde = 0.401
+ moin = 15.773 cgsl = {9.82591E-12/sw_func_tox_hv_ratio} cgdl = {9.82591E-12/sw_func_tox_hv_ratio}
+ ijthsrev = 0.1 ijthsfwd = 0.1 xjbvs = 1
+ bvs = 12.69 jss = 2.1483E-5 jsws = 4.02E-12
+ cjs = {sw_psd_nw_cj} mjs = 0.33956 mjsws = 0.24676
+ cjsws = {9.960545E-11*sw_func_psd_nw_cj} cjswgs = {1.47314E-10*sw_func_psd_nw_cj} mjswgs = 0.81
+ pbs = 0.6587 pbsws = 1 pbswgs = 3
+ xrcrg1 = 12 xrcrg2 = 1 rbpb = 50
+ rbpd = 50 rbps = 50 rbdb = 50
+ rbsb = 50 gbmin = 1E-12 tnom = 30
+ ute = -1.273991 lute = -1.698563E-7 wute = -4.933512E-7
+ pute = 4.485796E-13 kt1 = -0.491697 lkt1 = -1.257524E-7
+ wkt1 = -9.906651E-8 pkt1 = 9.007622E-14 kt1l = 0
+ kt2 = -0.019032 ua1 = 5.524E-10 ub1 = -3.075962E-18
+ lub1 = -4.682071E-25 wub1 = -4.548143E-24 pub1 = 4.135399E-30
+ uc1 = -1.092E-10 at = 2.309122E5 lat = -0.182679
+ wat = 0.207346 pat = -1.885295E-7 prt = 0
+ njs = 1.3632 xtis = 10 tpb = 1.671E-3
+ tpbsw = 0 tpbswg = 0 tcj = 9.6E-4
+ tcjsw = 3E-5 tcjswg = 0 tvoff = 0
+ tvfbsdoff = 0 saref = 3E-6 sbref = 3E-6
+ wlod = 0 ku0 = 7E-8 kvsat = 0.4
+ kvth0 = 3.5E-8 tku0 = 0 llodku0 = 0
+ wlodku0 = 1 llodvth = 0 wlodvth = 1
+ lku0 = 0 wku0 = 0 pku0 = 0
+ lkvth0 = 0 wkvth0 = 6.5E-7 pkvth0 = 0
+ stk2 = 0 lodk2 = 1 steta0 = 0
+ lodeta0 = 1

.model phv_model.26 pmos
+ level = 54 lmin = 8E-7 lmax = 1E-6 wmin = 3E-6
+ wmax = 7E-6 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 1.175E-8
+ toxm = 1.175E-8 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 1E23 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {1.2277E-8+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {4.5375E-8-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = -4.7338E-9 dwb = 0 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = -1.043407 lvth0 = 4.173358E-8
+ wvth0 = 2.555533E-7 pvth0 = -1.24176E-13 k1 = 0.598314
+ lk1 = -1.720624E-8 wk1 = -5.630602E-8 pk1 = 5.119625E-14
+ k2 = 1.32716E-2 lk2 = 1.859511E-8 wk2 = 5.590807E-8
+ pk2 = -5.532876E-14 k3 = -2.2405 k3b = -0.172
+ w0 = 0 lpe0 = 0 lpeb = 0
+ vbm = -3 dvtp0 = 0 dvtp1 = 0
+ dvt0 = 4.657 dvt1 = 0.34864 dvt2 = -0.030206
+ dvt0w = -2.2 dvt1w = 1.0163E6 dvt2w = 0
+ vfbsdoff = 0 u0 = 1.24541E-2 lu0 = 5.828756E-9
+ wu0 = 1.399017E-8 pu0 = -1.734315E-14 ua = -2.668779E-9
+ lua = 3.926832E-15 wua = 1.284637E-14 pua = -1.168408E-20
+ ub = 6.056562E-18 lub = -4.838328E-24 wub = -1.614576E-23
+ pub = 1.439618E-29 uc = 1.104288E-11 luc = -1.057307E-17
+ wuc = -3.45995E-17 puc = 3.145959E-23 ud = 0
+ up = 0 lp = 1 eu = 1.67
+ vsat = -2.103171E4 lvsat = 6.26662E-2 wvsat = 0.20507
+ pvsat = -1.864598E-7 a0 = 0.691766 la0 = 1.06122E-7
+ wa0 = 4.599777E-7 pa0 = -3.157604E-13 ags = 0.771528
+ lags = -2.595556E-8 wags = -2.052333E-7 pags = 7.722938E-14
+ b0 = 0 b1 = 0 keta = -0.205152
+ lketa = 1.095464E-7 wketa = 3.584817E-7 pketa = -3.259495E-13
+ a1 = 0 a2 = 0.5 rdsw = 788.47
+ rdswmin = 0 rdw = 0 rdwmin = 0
+ rsw = 0 rswmin = 0 prwb = 0.053538
+ prwg = 0 wr = 1 voff = -0.108271
+ lvoff = 2.77462E-8 wvoff = 9.079718E-8 pvoff = -8.255733E-14
+ voffl = 0 minv = 0 nfactor = 1.662337
+ lnfactor = 5.904103E-9 wnfactor = 3.675495E-8 pnfactor = -1.756734E-14
+ eta0 = -6.54543E-3 leta0 = 8.32591E-11 weta0 = 4.558481E-8
+ peta0 = -2.47733E-16 etab = 1.315806E-3 letab = -1.196396E-9
+ wetab = -3.915109E-9 petab = 3.559812E-15 dsub = 2.392177
+ ldsub = -1.514487E-6 wdsub = -6.228166E-6 pdsub = 4.506274E-12
+ cit = -2.592084E-5 lcit = 2.811478E-11 wcit = 9.20033E-11
+ pcit = -8.3654E-17 cdsc = 0 cdscb = 0
+ cdscd = 0 pclm = 2.631067 lpclm = -1.298368E-6
+ wpclm = -4.248802E-6 ppclm = 3.863223E-12 pdiblc1 = 0.044364
+ lpdiblc1 = 3.229315E-7 wpdiblc1 = 1.056767E-6 ppdiblc1 = -9.608651E-13
+ pdiblc2 = -5.97464E-2 lpdiblc2 = 5.569392E-8 wpdiblc2 = 1.822538E-7
+ ppdiblc2 = -1.657143E-13 pdiblcb = -0.025 drout = 0.280167
+ ldrout = 1.186778E-7 wdrout = 3.883632E-7 pdrout = -3.531193E-13
+ pscbe1 = -3.221505E8 lpscbe1 = 565.217802 wpscbe1 = 1.849629E3
+ ppscbe1 = -1.681775E-3 pscbe2 = 2.105385E-8 lpscbe2 = -5.909468E-15
+ wpscbe2 = -1.933825E-14 ppscbe2 = 1.75833E-20 pvag = 0
+ delta = 0.01 fprout = 0 pdits = 0
+ pditsl = 0 pditsd = 0 lambda = 0
+ vtl = 0 lc = 5E-9 xn = 3
+ alpha0 = 3.805651E-4 lalpha0 = -2.843697E-10 walpha0 = -9.305764E-10
+ palpha0 = 8.461266E-16 alpha1 = 0 beta0 = 79.875246
+ lbeta0 = -2.702502E-5 wbeta0 = -8.843716E-5 pbeta0 = 8.041149E-11
+ aigbacc = 0.43 bigbacc = 0.054 cigbacc = 0.075
+ nigbacc = 1 aigbinv = 0.35 bigbinv = 0.03
+ cigbinv = 6E-3 eigbinv = 1.1 nigbinv = 3
+ aigc = 0.43 bigc = 0.054 cigc = 0.075
+ aigsd = 0.43 bigsd = 0.054 cigsd = 0.075
+ dlcig = 0 nigc = 1 poxedge = 1
+ pigcd = 1 ntox = 1 toxref = 1.175E-8
+ agidl = -8.555526E-9 lagidl = 1.694534E-14 wagidl = 4.335203E-14
+ pagidl = -5.041994E-20 bgidl = 1.049751E9 lbgidl = 665.757934
+ wbgidl = 1.529524E3 pbgidl = -1.980927E-3 cgidl = -982.605212
+ lcgidl = 8.546892E-4 wcgidl = 5.661099E-3 pcgidl = -2.543082E-9
+ egidl = 2.621504 legidl = -1.675316E-6 wegidl = -5.482333E-6
+ pegidl = 4.984811E-12 noia = 3E40 noib = 8.53E24
+ noic = 8.4E7 em = 4.1E7 af = 1
+ ef = 0.88 kf = 0 lintnoi = 0
+ tnoia = 1.5 tnoib = 3.5 ntnoi = 1
+ rnoia = 0.577 rnoib = 0.37 xpart = 0
+ cgso = {1.94171E-10/sw_func_tox_hv_ratio} cgdo = {1.94171E-10/sw_func_tox_hv_ratio} cgbo = {0/sw_func_tox_hv_ratio}
+ ckappas = 0.6 cf = 1.2E-11 clc = 1E-7
+ cle = 0.6 dlc = 4.4983E-8 dwc = 0
+ vfbcv = -0.144689 noff = 4 voffcv = 0
+ acde = 0.401 moin = 15.773 cgsl = {9.82591E-12/sw_func_tox_hv_ratio}
+ cgdl = {9.82591E-12/sw_func_tox_hv_ratio} ijthsrev = 0.1 ijthsfwd = 0.1
+ xjbvs = 1 bvs = 12.69 jss = 2.1483E-5
+ jsws = 4.02E-12 cjs = {sw_psd_nw_cj} mjs = 0.33956
+ mjsws = 0.24676 cjsws = {9.960545E-11*sw_func_psd_nw_cj} cjswgs = {1.47314E-10*sw_func_psd_nw_cj}
+ mjswgs = 0.81 pbs = 0.6587 pbsws = 1
+ pbswgs = 3 xrcrg1 = 12 xrcrg2 = 1
+ rbpb = 50 rbpd = 50 rbps = 50
+ rbdb = 50 rbsb = 50 gbmin = 1E-12
+ tnom = 30 ute = -1.343301 lute = -1.068362E-7
+ wute = -3.496125E-7 pute = 3.178852E-13 kt1 = -0.546514
+ lkt1 = -7.59099E-8 wkt1 = -2.484089E-7 pkt1 = 2.258658E-13
+ kt1l = 0 kt2 = -0.019032 ua1 = 5.524E-10
+ ub1 = -3.5909E-18 uc1 = -1.092E-10 at = 6.092084E4
+ lat = -2.81148E-2 wat = -9.20033E-2 pat = 8.3654E-8
+ prt = 0 njs = 1.3632 xtis = 10
+ tpb = 1.671E-3 tpbsw = 0 tpbswg = 0
+ tcj = 9.6E-4 tcjsw = 3E-5 tcjswg = 0
+ tvoff = 0 tvfbsdoff = 0 saref = 2.81E-6
+ sbref = 2.81E-6 wlod = 0 ku0 = 7E-8
+ kvsat = 0.4 kvth0 = 3.5E-8 tku0 = 0
+ llodku0 = 0 wlodku0 = 1 llodvth = 0
+ wlodvth = 1 lku0 = 0 wku0 = 0
+ pku0 = 0 lkvth0 = 0 wkvth0 = 6.5E-7
+ pkvth0 = 0 stk2 = 0 lodk2 = 1
+ steta0 = 0 lodeta0 = 1

.model phv_model.27 pmos
+ level = 54 lmin = 6E-7 lmax = 8E-7 wmin = 3E-6
+ wmax = 7E-6 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 1.175E-8
+ toxm = 1.175E-8 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 1E23 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {1.2277E-8+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {4.5375E-8-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = -4.7338E-9 dwb = 0 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = -0.965066 lvth0 = -1.382989E-8
+ wvth0 = -5.554389E-8 pvth0 = 9.646967E-14 k1 = 0.568258
+ lk1 = 4.110682E-9 wk1 = 5.630602E-8 pk1 = -2.867384E-14
+ k2 = 5.48686E-2 lk2 = -1.090757E-8 wk2 = -1.293777E-7
+ pk2 = 7.608518E-14 k3 = -2.2405 k3b = -0.172
+ w0 = 0 lpe0 = 0 lpeb = 0
+ vbm = -3 dvtp0 = 0 dvtp1 = 0
+ dvt0 = 4.657 dvt1 = 0.34864 dvt2 = -0.030206
+ dvt0w = -2.2 dvt1w = 1.0163E6 dvt2w = 0
+ vfbsdoff = 0 u0 = 2.14171E-2 lu0 = -5.282092E-10
+ wu0 = -1.565754E-8 pu0 = 3.684495E-15 ua = 4.185805E-9
+ lua = -9.347815E-16 wua = -1.282102E-14 pua = 6.520518E-21
+ ub = -2.603941E-18 lub = 1.304134E-24 wub = 1.697811E-23
+ pub = -9.096917E-30 uc = -7.425984E-12 luc = 2.525974E-18
+ wuc = 3.45995E-17 puc = -1.761979E-23 ud = 0
+ up = 0 lp = 1 eu = 1.67
+ vsat = 1.161687E5 lvsat = -3.46432E-2 wvsat = -0.398542
+ pvsat = 2.416521E-7 a0 = 0.835999 la0 = 3.825084E-9
+ wa0 = 5.239404E-8 pa0 = -2.668167E-14 ags = 0.770101
+ lags = -2.494339E-8 wags = -3.416618E-7 pags = 1.739913E-13
+ b0 = 0 b1 = 0 keta = 2.81837E-2
+ lketa = -5.594692E-8 wketa = -6.513233E-7 pketa = 3.902547E-13
+ a1 = 0 a2 = 0.5 rdsw = 788.47
+ rdswmin = 0 rdw = 0 rdwmin = 0
+ rsw = 0 rswmin = 0 prwb = 0.053538
+ prwg = 0 wr = 1 voff = -5.98046E-2
+ lvoff = -6.628746E-9 wvoff = -9.079718E-8 pvoff = 4.623846E-14
+ voffl = 0 minv = 0 nfactor = 1.840578
+ lnfactor = -1.205128E-7 wnfactor = -1.173253E-6 pnfactor = 8.406308E-13
+ eta0 = -0.02259 leta0 = 1.146285E-8 weta0 = 1.579722E-7
+ peta0 = -7.995851E-14 etab = -3.710414E-4 wetab = 1.104014E-9
+ dsub = 0.211063 ldsub = 3.246834E-8 wdsub = 4.447348E-7
+ pdsub = -2.264812E-13 cit = 2.318959E-5 lcit = -6.716801E-12
+ wcit = -9.20033E-11 pcit = 4.685268E-17 cdsc = 0
+ cdscb = 0 cdscd = 0 pclm = 0.363104
+ lpclm = 3.101852E-7 wpclm = 4.248771E-6 ppclm = -2.16368E-12
+ pdiblc1 = 0.608455 lpdiblc1 = -7.71504E-8 wpdiblc1 = -1.056767E-6
+ ppdiblc1 = 5.381584E-13 pdiblc2 = 3.75388E-2 lpdiblc2 = -1.330563E-8
+ wpdiblc2 = -1.822538E-7 ppdiblc2 = 9.281274E-14 pdiblcb = -0.025
+ drout = 0.487471 ldrout = -2.835288E-8 wdrout = -3.883632E-7
+ pdrout = 1.97774E-13 pscbe1 = 6.651628E8 lpscbe1 = -135.034161
+ wpscbe1 = -1.849629E3 ppscbe1 = 9.419235E-4 pscbe2 = 1.073128E-8
+ lpscbe2 = 1.41181E-15 wpscbe2 = 1.933825E-14 ppscbe2 = -9.848003E-21
+ pvag = 0 delta = 0.01 fprout = 0
+ pdits = 0 pditsl = 0 pditsd = 0
+ lambda = 0 vtl = 0 lc = 5E-9
+ xn = 3 alpha0 = -1.161673E-4 lalpha0 = 6.793774E-11
+ walpha0 = 9.305764E-10 palpha0 = -4.73896E-16 alpha1 = 0
+ beta0 = 32.668378 lbeta0 = 6.456451E-6 wbeta0 = 8.843716E-5
+ pbeta0 = -4.503662E-11 aigbacc = 0.43 bigbacc = 0.054
+ cigbacc = 0.075 nigbacc = 1 aigbinv = 0.35
+ bigbinv = 0.03 cigbinv = 6E-3 eigbinv = 1.1
+ nigbinv = 3 aigc = 0.43 bigc = 0.054
+ cigc = 0.075 aigsd = 0.43 bigsd = 0.054
+ cigsd = 0.075 dlcig = 0 nigc = 1
+ poxedge = 1 pigcd = 1 ntox = 1
+ toxref = 1.175E-8 agidl = 2.609387E-8 lagidl = -7.629748E-15
+ wagidl = -1.027753E-13 pagidl = 5.32209E-20 bgidl = 2.449633E9
+ lbgidl = -327.108202 wbgidl = -4.480561E3 pbgidl = 2.281726E-3
+ cgidl = -535.167538 lcgidl = 5.373441E-4 wcgidl = 7.360264E-3
+ pcgidl = -3.748215E-9 egidl = -0.30491 legidl = 4.002437E-7
+ wegidl = 5.482333E-6 pegidl = -2.791878E-12 noia = 3E40
+ noib = 8.53E24 noic = 8.4E7 em = 4.1E7
+ af = 1 ef = 0.88 kf = 0
+ lintnoi = 0 tnoia = 1.5 tnoib = 3.5
+ ntnoi = 1 rnoia = 0.577 rnoib = 0.37
+ xpart = 0 cgso = {1.94171E-10/sw_func_tox_hv_ratio} cgdo = {1.94171E-10/sw_func_tox_hv_ratio}
+ cgbo = {0/sw_func_tox_hv_ratio} ckappas = 0.6 cf = 1.2E-11
+ clc = 1E-7 cle = 0.6 dlc = 4.4983E-8
+ dwc = 0 vfbcv = -0.144689 noff = 4
+ voffcv = 0 acde = 0.401 moin = 15.773
+ cgsl = {9.82591E-12/sw_func_tox_hv_ratio} cgdl = {9.82591E-12/sw_func_tox_hv_ratio} ijthsrev = 0.1
+ ijthsfwd = 0.1 xjbvs = 1 bvs = 12.69
+ jss = 2.1483E-5 jsws = 4.02E-12 cjs = {sw_psd_nw_cj}
+ mjs = 0.33956 mjsws = 0.24676 cjsws = {9.960545E-11*sw_func_psd_nw_cj}
+ cjswgs = {1.47314E-10*sw_func_psd_nw_cj} mjswgs = 0.81 pbs = 0.6587
+ pbsws = 1 pbswgs = 3 xrcrg1 = 12
+ xrcrg2 = 1 rbpb = 50 rbpd = 50
+ rbps = 50 rbdb = 50 rbsb = 50
+ gbmin = 1E-12 tnom = 30 ute = -1.487304
+ lute = -4.701761E-9 wute = 5.234492E-8 pute = 3.279688E-14
+ kt1 = -0.682862 lkt1 = 2.079522E-8 wkt1 = 2.745685E-7
+ pkt1 = -1.450559E-13 kt1l = 0 kt2 = -0.019032
+ ua1 = 5.524E-10 ub1 = -3.038403E-18 lub1 = -3.918582E-25
+ wub1 = -3.85391E-24 pub1 = 2.733385E-30 uc1 = 1.903526E-11
+ luc1 = -9.095086E-17 wuc1 = -8.944981E-16 puc1 = 6.344228E-22
+ at = -1.447996E3 lat = 1.61203E-2 wat = 0.184487
+ pat = -1.124464E-7 prt = 0 njs = 1.3632
+ xtis = 10 tpb = 1.671E-3 tpbsw = 0
+ tpbswg = 0 tcj = 9.6E-4 tcjsw = 3E-5
+ tcjswg = 0 tvoff = 0 tvfbsdoff = 0
+ saref = 2.81E-6 sbref = 2.81E-6 wlod = 0
+ ku0 = 7E-8 kvsat = 0.4 kvth0 = 3.5E-8
+ tku0 = 0 llodku0 = 0 wlodku0 = 1
+ llodvth = 0 wlodvth = 1 lku0 = 0
+ wku0 = 0 pku0 = 0 lkvth0 = 0
+ wkvth0 = 6.5E-7 pkvth0 = 0 stk2 = 0
+ lodk2 = 1 steta0 = 0 lodeta0 = 1

.model phv_model.28 pmos
+ level = 54 lmin = 5E-7 lmax = 6E-7 wmin = 3E-6
+ wmax = 7E-6 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 1.175E-8
+ toxm = 1.175E-8 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 1E23 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {1.2277E-8+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {4.5375E-8-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = -4.7338E-9 dwb = 0 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = -0.924231 lvth0 = -3.462519E-8
+ wvth0 = 5.237022E-7 pvth0 = -1.985114E-13 k1 = 0.398285
+ lk1 = 9.066931E-8 wk1 = 6.221862E-7 pk1 = -3.168483E-13
+ k2 = 2.40833E-2 lk2 = 4.769858E-9 wk2 = 1.33396E-8
+ pk2 = 3.40639E-15 k3 = -2.2405 k3b = -0.172
+ w0 = 0 lpe0 = 0 lpeb = 0
+ vbm = -3 dvtp0 = 0 dvtp1 = 0
+ dvt0 = 4.657 dvt1 = 0.34864 dvt2 = -0.030206
+ dvt0w = -2.2 dvt1w = 1.0163E6 dvt2w = 0
+ vfbsdoff = 0 u0 = 2.48403E-2 lu0 = -2.271509E-9
+ wu0 = -5.082386E-8 pu0 = 2.159294E-14 ua = 4.479128E-9
+ lua = -1.084156E-15 wua = -9.511943E-15 pua = 4.835371E-21
+ ub = -2.451637E-18 lub = 1.226573E-24 wub = -8.916258E-25
+ pub = 3.244181E-33 uc = -8.445744E-11 luc = 4.175424E-17
+ wuc = 6.523081E-16 puc = -3.321879E-22 ud = 0
+ up = 0 lp = 1 eu = 1.67
+ vsat = 1.718738E5 lvsat = -0.063011 wvsat = -0.898857
+ pvsat = 4.964375E-7 a0 = 0.265109 la0 = 2.945509E-7
+ wa0 = 7.194426E-7 pa0 = -3.663761E-13 ags = -4.67023
+ lags = 2.745545E-6 wags = 2.250913E-5 pags = -1.146277E-11
+ b0 = 0 b1 = 0 keta = 0.194146
+ lketa = -1.404634E-7 wketa = -1.218635E-6 pketa = 6.79158E-13
+ a1 = 0 a2 = 0.5 rdsw = 788.47
+ rdswmin = 0 rdw = 0 rdwmin = 0
+ rsw = 0 rswmin = 0 prwb = 0.053538
+ prwg = 0 wr = 1 voff = -1.27682E-2
+ lvoff = -3.058208E-8 wvoff = 4.008423E-7 pvoff = -2.041289E-13
+ voffl = 0 minv = 0 nfactor = 0.395692
+ lnfactor = 6.152949E-7 wnfactor = 5.953133E-6 pnfactor = -2.788481E-12
+ eta0 = -0.13398 leta0 = 6.818827E-8 weta0 = -1.348738E-6
+ peta0 = 6.873337E-13 etab = -2.04035E-2 letab = 1.020151E-8
+ wetab = 2.446797E-7 petab = -1.240409E-13 dsub = 0.296008
+ ldsub = -1.078994E-8 wdsub = -2.862481E-7 pdsub = 1.457719E-13
+ cit = 4.568377E-5 lcit = -1.817196E-11 wcit = -1.061751E-10
+ pcit = 5.406968E-17 cdsc = 0 cdscb = 0
+ cdscd = 0 pclm = -2.744381 lpclm = 1.892672E-6
+ wpclm = 1.552163E-5 ppclm = -7.904386E-12 pdiblc1 = 0.80501
+ lpdiblc1 = -1.772456E-7 wpdiblc1 = 2.223259E-6 ppdiblc1 = -1.132195E-12
+ pdiblc2 = 3.55024E-2 lpdiblc2 = -1.22686E-8 wpdiblc2 = 2.064797E-8
+ ppdiblc2 = -1.051498E-14 pdiblcb = -0.633851 lpdiblcb = 3.100572E-7
+ wpdiblcb = 4.247005E-6 ppdiblcb = -2.162787E-12 drout = -1.177085
+ ldrout = 8.193221E-7 wdrout = -2.1319E-6 pdrout = 1.08567E-12
+ pscbe1 = 5.702684E8 lpscbe1 = -86.709162 wpscbe1 = -121.180211
+ ppscbe1 = 6.171102E-5 pscbe2 = 9.651958E-9 lpscbe2 = 1.961456E-15
+ wpscbe2 = -1.197974E-15 ppscbe2 = 6.100682E-22 pvag = 0
+ delta = 0.01 fprout = 0 pdits = 0
+ pditsl = 0 pditsd = 0 lambda = 0
+ vtl = 0 lc = 5E-9 xn = 3
+ alpha0 = -6.054351E-4 lalpha0 = 3.170974E-10 walpha0 = 2.062669E-9
+ palpha0 = -1.050414E-15 alpha1 = 3.044253E-10 lalpha1 = -1.550286E-16
+ walpha1 = -2.123502E-15 palpha1 = 1.081394E-21 beta0 = -150.208876
+ lbeta0 = 9.958669E-5 wbeta0 = 1.097522E-3 pbeta0 = -5.58913E-10
+ aigbacc = 0.43 bigbacc = 0.054 cigbacc = 0.075
+ nigbacc = 1 aigbinv = 0.35 bigbinv = 0.03
+ cigbinv = 6E-3 eigbinv = 1.1 nigbinv = 3
+ aigc = 0.43 bigc = 0.054 cigc = 0.075
+ aigsd = 0.43 bigsd = 0.054 cigsd = 0.075
+ dlcig = 0 nigc = 1 poxedge = 1
+ pigcd = 1 ntox = 1 toxref = 1.175E-8
+ agidl = 3.341201E-8 lagidl = -1.135651E-14 wagidl = -1.207081E-13
+ pagidl = 6.235315E-20 bgidl = 1.804617E9 lbgidl = 1.366572
+ wbgidl = 7.158326E3 pbgidl = -3.645378E-3 cgidl = 3.74557E3
+ lcgidl = -1.642622E-3 wcgidl = -1.26225E-2 pcgidl = 6.42802E-9
+ egidl = 3.790328 legidl = -1.685257E-6 wegidl = -2.834305E-5
+ pegidl = 1.44337E-11 noia = 3E40 noib = 8.53E24
+ noic = 8.4E7 em = 4.1E7 af = 1
+ ef = 0.88 kf = 0 lintnoi = 0
+ tnoia = 1.5 tnoib = 3.5 ntnoi = 1
+ rnoia = 0.577 rnoib = 0.37 xpart = 0
+ cgso = {1.94171E-10/sw_func_tox_hv_ratio} cgdo = {1.94171E-10/sw_func_tox_hv_ratio} cgbo = {0/sw_func_tox_hv_ratio}
+ ckappas = 0.6 cf = 1.2E-11 clc = 1E-7
+ cle = 0.6 dlc = 4.4983E-8 dwc = 0
+ vfbcv = -0.144689 noff = 4 voffcv = 0
+ acde = 0.401 moin = 15.773 cgsl = {9.82591E-12/sw_func_tox_hv_ratio}
+ cgdl = {9.82591E-12/sw_func_tox_hv_ratio} ijthsrev = 0.1 ijthsfwd = 0.1
+ xjbvs = 1 bvs = 12.69 jss = 2.1483E-5
+ jsws = 4.02E-12 cjs = {sw_psd_nw_cj} mjs = 0.33956
+ mjsws = 0.24676 cjsws = {9.960545E-11*sw_func_psd_nw_cj} cjswgs = {1.47314E-10*sw_func_psd_nw_cj}
+ mjswgs = 0.81 pbs = 0.6587 pbsws = 1
+ pbswgs = 3 xrcrg1 = 12 xrcrg2 = 1
+ rbpb = 50 rbpd = 50 rbps = 50
+ rbdb = 50 rbsb = 50 gbmin = 1E-12
+ tnom = 30 ute = -1.700142 lute = 1.036858E-7
+ wute = -1.528967E-6 pute = 8.3808E-13 kt1 = -0.757162
+ lkt1 = 5.863234E-8 wkt1 = -3.496094E-7 pkt1 = 1.728067E-13
+ kt1l = 0 kt2 = -0.019032 ua1 = 5.52E-10
+ ub1 = -1.278633E-17 lub1 = 4.572275E-24 wub1 = 2.329433E-23
+ pub1 = -1.109185E-29 uc1 = -6.427491E-10 luc1 = 2.460628E-16
+ wuc1 = 1.788996E-15 puc1 = -7.321467E-22 at = 8.01643E4
+ lat = -2.54407E-2 wat = -0.184967 pat = 7.569755E-8
+ prt = 0 njs = 1.3632 xtis = 10
+ tpb = 1.671E-3 tpbsw = 0 tpbswg = 0
+ tcj = 9.6E-4 tcjsw = 3E-5 tcjswg = 0
+ tvoff = 0 tvfbsdoff = 0 saref = 2.02E-6
+ sbref = 2.01E-6 wlod = 0 ku0 = 7E-8
+ kvsat = 0.4 kvth0 = 3.5E-8 tku0 = 0
+ llodku0 = 0 wlodku0 = 1 llodvth = 0
+ wlodvth = 1 lku0 = 0 wku0 = 0
+ pku0 = 0 lkvth0 = 0 wkvth0 = 6.5E-7
+ pkvth0 = 0 stk2 = 0 lodk2 = 1
+ steta0 = 0 lodeta0 = 1

.model phv_model.29 pmos
+ level = 54 lmin = 8E-6 lmax = 2.02E-5 wmin = 1E-6
+ wmax = 3E-6 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 1.175E-8
+ toxm = 1.175E-8 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 1E23 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {1.2277E-8+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {4.5375E-8-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = -4.7338E-9 dwb = 0 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = -0.997895 wvth0 = 3.678035E-8
+ k1 = 0.600263 wk1 = -1.503436E-8 k2 = 2.48199E-2
+ wk2 = 3.994424E-10 k3 = -2.2405 k3b = -0.172
+ w0 = 0 lpe0 = 0 lpeb = 0
+ vbm = -3 dvtp0 = 0 dvtp1 = 0
+ dvt0 = 4.657 dvt1 = 0.34864 dvt2 = -0.030206
+ dvt0w = -2.2 dvt1w = 1.0163E6 dvt2w = 0
+ vfbsdoff = 0 u0 = 2.03215E-2 wu0 = -1.676694E-9
+ ua = 2.840714E-9 wua = -5.75742E-16 ub = -4.165952E-19
+ wub = 6.479187E-25 uc = -3.746677E-11 wuc = -7.454174E-18
+ ud = 0 up = 0 lp = 1
+ eu = 1.67 vsat = 2.584507E5 wvsat = -0.173917
+ a0 = 1.252938 wa0 = -3.380042E-7 ags = 0.169981
+ wags = -3.158903E-8 b0 = 0 b1 = 0
+ keta = -7.801043E-3 wketa = -3.715055E-10 a1 = 0
+ a2 = 0.5 rdsw = 788.47 rdswmin = 0
+ rdw = 0 rdwmin = 0 rsw = 0
+ rswmin = 0 prwb = 0.053538 prwg = 0
+ wr = 1 voff = -8.61446E-2 wvoff = -2.100671E-8
+ voffl = 0 minv = 0 nfactor = 1.808434
+ wnfactor = -2.046618E-7 eta0 = 0.08 etab = -0.07
+ dsub = 0.56 cit = 1.243862E-5 wcit = -7.255967E-12
+ cdsc = 0 cdscb = 0 cdscd = 0
+ pclm = 8.35312E-2 pdiblc1 = 0.39 pdiblc2 = 2.698253E-3
+ wpdiblc2 = 7.216479E-10 pdiblcb = -0.025 drout = 0.56
+ pscbe1 = 3.868723E8 wpscbe1 = -158.173149 pscbe2 = 1.499872E-8
+ pvag = 0 delta = 0.01 fprout = 0
+ pdits = 0 pditsl = 0 pditsd = 0
+ lambda = 0 vtl = 0 lc = 5E-9
+ xn = 3 alpha0 = 4.404613E-5 walpha0 = 1.970061E-11
+ alpha1 = 0 beta0 = 37.888825 wbeta0 = 1.122399E-6
+ aigbacc = 0.43 bigbacc = 0.054 cigbacc = 0.075
+ nigbacc = 1 aigbinv = 0.35 bigbinv = 0.03
+ cigbinv = 6E-3 eigbinv = 1.1 nigbinv = 3
+ aigc = 0.43 bigc = 0.054 cigc = 0.075
+ aigsd = 0.43 bigsd = 0.054 cigsd = 0.075
+ dlcig = 0 nigc = 1 poxedge = 1
+ pigcd = 1 ntox = 1 toxref = 1.175E-8
+ agidl = 1.222665E-8 wagidl = 7.582486E-15 bgidl = 1.900216E9
+ wbgidl = -370.489688 cgidl = 804.9108 wcgidl = 5.804774E-4
+ egidl = 0.290441 wegidl = 1.199305E-6 noia = 3E40
+ noib = 8.53E24 noic = 8.4E7 em = 4.1E7
+ af = 1 ef = 0.88 kf = 0
+ lintnoi = 0 tnoia = 1.5 tnoib = 3.5
+ ntnoi = 1 rnoia = 0.577 rnoib = 0.37
+ xpart = 0 cgso = {1.94171E-10/sw_func_tox_hv_ratio} cgdo = {1.94171E-10/sw_func_tox_hv_ratio}
+ cgbo = {0/sw_func_tox_hv_ratio} ckappas = 0.6 cf = 1.2E-11
+ clc = 1E-7 cle = 0.6 dlc = 4.4983E-8
+ dwc = 0 vfbcv = -0.144689 noff = 4
+ voffcv = 0 acde = 0.401 moin = 15.773
+ cgsl = {9.82591E-12/sw_func_tox_hv_ratio} cgdl = {9.82591E-12/sw_func_tox_hv_ratio} ijthsrev = 0.1
+ ijthsfwd = 0.1 xjbvs = 1 bvs = 12.69
+ jss = 2.1483E-5 jsws = 4.02E-12 cjs = {sw_psd_nw_cj}
+ mjs = 0.33956 mjsws = 0.24676 cjsws = {9.960545E-11*sw_func_psd_nw_cj}
+ cjswgs = {1.47314E-10*sw_func_psd_nw_cj} mjswgs = 0.81 pbs = 0.6587
+ pbsws = 1 pbswgs = 3 xrcrg1 = 12
+ xrcrg2 = 1 rbpb = 50 rbpd = 50
+ rbps = 50 rbdb = 50 rbsb = 50
+ gbmin = 1E-12 tnom = 30 ute = -1.526346
+ wute = -2.902387E-8 kt1 = -0.585754 wkt1 = 2.902387E-8
+ kt1l = 0 kt2 = -0.019032 ua1 = 2.2096E-11
+ ub1 = -3.948506E-18 wub1 = 8.503994E-25 uc1 = -1.092E-10
+ at = 5.94E5 wat = -0.432035 prt = 0
+ njs = 1.3632 xtis = 10 tpb = 1.671E-3
+ tpbsw = 0 tpbswg = 0 tcj = 9.6E-4
+ tcjsw = 3E-5 tcjswg = 0 tvoff = 0
+ tvfbsdoff = 0 saref = 3E-6 sbref = 3E-6
+ wlod = 0 ku0 = 7E-8 kvsat = 0.4
+ kvth0 = 3.5E-8 tku0 = 0 llodku0 = 0
+ wlodku0 = 1 llodvth = 0 wlodvth = 1
+ lku0 = 0 wku0 = 0 pku0 = 0
+ lkvth0 = 0 wkvth0 = 6.5E-7 pkvth0 = 0
+ stk2 = 0 lodk2 = 1 steta0 = 0
+ lodeta0 = 1

.model phv_model.30 pmos
+ level = 54 lmin = 4E-6 lmax = 8E-6 wmin = 1E-6
+ wmax = 3E-6 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 1.175E-8
+ toxm = 1.175E-8 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 1E23 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {1.2277E-8+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {4.5375E-8-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = -4.7338E-9 dwb = 0 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = -0.99492 lvth0 = -2.353109E-8
+ wvth0 = 2.049181E-8 pvth0 = 1.288301E-13 k1 = 0.623219
+ lk1 = -1.815659E-7 wk1 = -5.673149E-8 pk1 = 3.29793E-13
+ k2 = 1.98284E-2 lk2 = 3.947872E-8 wk2 = 1.132875E-8
+ pk2 = -8.64426E-14 k3 = -2.2405 k3b = -0.172
+ w0 = 0 lpe0 = 0 lpeb = 0
+ vbm = -3 dvtp0 = 0 dvtp1 = 0
+ dvt0 = 4.657 dvt1 = 0.34864 dvt2 = -0.030206
+ dvt0w = -2.2 dvt1w = 1.0163E6 dvt2w = 0
+ vfbsdoff = 0 u0 = 1.87624E-2 lu0 = 1.233116E-8
+ wu0 = 5.629233E-10 pu0 = -1.77137E-14 ua = 2.244397E-9
+ lua = 4.716418E-15 wua = 2.764605E-16 pua = -6.740282E-21
+ ub = 1.799087E-19 lub = -4.717898E-24 wub = -5.877238E-26
+ pub = 5.589396E-30 uc = -4.748145E-11 luc = 7.920863E-17
+ wuc = -1.2182E-17 puc = 3.739359E-23 ud = 0
+ up = 0 lp = 1 eu = 1.67
+ vsat = 3.867309E5 lvsat = -1.0146 wvsat = -0.33725
+ pvsat = 1.291846E-6 a0 = 1.614328 la0 = -2.858328E-6
+ wa0 = -6.534178E-7 pa0 = 2.494685E-12 ags = 0.183711
+ lags = -1.086002E-7 wags = -4.531548E-8 pags = 1.085659E-13
+ b0 = 0 b1 = 0 keta = -4.167981E-3
+ lketa = -2.87348E-8 wketa = -2.346871E-9 pketa = 1.562366E-14
+ a1 = 0 a2 = 0.5 rdsw = 788.47
+ rdswmin = 0 rdw = 0 rdwmin = 0
+ rsw = 0 rswmin = 0 prwb = 0.053538
+ prwg = 0 wr = 1 voff = -8.34259E-2
+ lvoff = -2.150317E-8 wvoff = -3.377304E-8 pvoff = 1.009721E-13
+ voffl = 0 minv = 0 nfactor = 1.828691
+ lnfactor = -1.602191E-7 wnfactor = -2.829361E-7 pnfactor = 6.19091E-13
+ eta0 = 0.08 etab = -0.07 dsub = 0.56
+ cit = 1.48219E-5 lcit = -1.885003E-11 wcit = -1.434731E-11
+ pcit = 5.608724E-17 cdsc = 0 cdscb = 0
+ cdscd = 0 pclm = -0.60959 lpclm = 5.482071E-6
+ wpclm = -1.152362E-7 ppclm = 9.114322E-13 pdiblc1 = 0.39
+ pdiblc2 = 4.074557E-3 lpdiblc2 = -1.088553E-8 wpdiblc2 = 1.426923E-9
+ ppdiblc2 = -5.5782E-15 pdiblcb = -0.025 drout = 0.56
+ pscbe1 = 7.268464E8 lpscbe1 = -2.68894E3 wpscbe1 = -490.124642
+ ppscbe1 = 2.625487E-3 pscbe2 = -3.009912E-8 lpscbe2 = 3.567164E-13
+ wpscbe2 = 4.398225E-14 ppscbe2 = -3.478923E-19 pvag = 0
+ delta = 0.01 fprout = 0 pdits = 0
+ pditsl = 0 pditsd = 0 lambda = 0
+ vtl = 0 lc = 5E-9 xn = 3
+ alpha0 = 5.431603E-5 lalpha0 = -8.122719E-11 walpha0 = 7.092629E-11
+ palpha0 = -4.051567E-16 alpha1 = 4.766578E-11 lalpha1 = -3.770006E-16
+ walpha1 = -1.418269E-16 palpha1 = 1.121745E-21 beta0 = 22.010958
+ lbeta0 = 1.25582E-4 wbeta0 = 5.09674E-5 pbeta0 = -3.942365E-10
+ aigbacc = 0.43 bigbacc = 0.054 cigbacc = 0.075
+ nigbacc = 1 aigbinv = 0.35 bigbinv = 0.03
+ cigbinv = 6E-3 eigbinv = 1.1 nigbinv = 3
+ aigc = 0.43 bigc = 0.054 cigc = 0.075
+ aigsd = 0.43 bigsd = 0.054 cigsd = 0.075
+ dlcig = 0 nigc = 1 poxedge = 1
+ pigcd = 1 ntox = 1 toxref = 1.175E-8
+ agidl = 2.652428E-8 lagidl = -1.130836E-13 wagidl = -1.932918E-14
+ pagidl = 2.128511E-19 bgidl = 1.752102E9 lbgidl = 1.171471E3
+ wbgidl = -180.157921 pbgidl = -1.505382E-3 cgidl = 866.455428
+ lcgidl = -4.867719E-4 wcgidl = 1.386054E-3 pcgidl = -6.37151E-9
+ egidl = 1.286651 legidl = -7.879273E-6 wegidl = -2.300968E-7
+ pegidl = 1.13055E-11 noia = 3E40 noib = 8.53E24
+ noic = 8.4E7 em = 4.1E7 af = 1
+ ef = 0.88 kf = 0 lintnoi = 0
+ tnoia = 1.5 tnoib = 3.5 ntnoi = 1
+ rnoia = 0.577 rnoib = 0.37 xpart = 0
+ cgso = {1.94171E-10/sw_func_tox_hv_ratio} cgdo = {1.94171E-10/sw_func_tox_hv_ratio} cgbo = {0/sw_func_tox_hv_ratio}
+ ckappas = 0.6 cf = 1.2E-11 clc = 1E-7
+ cle = 0.6 dlc = 4.4983E-8 dwc = 0
+ vfbcv = -0.144689 noff = 4 voffcv = 0
+ acde = 0.401 moin = 15.773 cgsl = {9.82591E-12/sw_func_tox_hv_ratio}
+ cgdl = {9.82591E-12/sw_func_tox_hv_ratio} ijthsrev = 0.1 ijthsfwd = 0.1
+ xjbvs = 1 bvs = 12.69 jss = 2.1483E-5
+ jsws = 4.02E-12 cjs = {sw_psd_nw_cj} mjs = 0.33956
+ mjsws = 0.24676 cjsws = {9.960545E-11*sw_func_psd_nw_cj} cjswgs = {1.47314E-10*sw_func_psd_nw_cj}
+ mjswgs = 0.81 pbs = 0.6587 pbsws = 1
+ pbswgs = 3 xrcrg1 = 12 xrcrg2 = 1
+ rbpb = 50 rbpd = 50 rbps = 50
+ rbdb = 50 rbsb = 50 gbmin = 1E-12
+ tnom = 30 ute = -1.427817 lute = -7.792861E-7
+ wute = -2.640311E-7 pute = 1.858731E-12 kt1 = -0.595288
+ lkt1 = 7.540011E-8 wkt1 = 5.738926E-8 pkt1 = -2.24349E-13
+ kt1l = 0 kt2 = -0.019032 ua1 = 2.2096E-11
+ ub1 = -3.49369E-18 lub1 = -3.59725E-24 wub1 = -2.38548E-25
+ pub1 = 8.612757E-30 uc1 = -1.092E-10 at = 9.453027E5
+ lat = -2.778541 wat = -0.840071 pat = 3.22726E-6
+ prt = 0 njs = 1.3632 xtis = 10
+ tpb = 1.671E-3 tpbsw = 0 tpbswg = 0
+ tcj = 9.6E-4 tcjsw = 3E-5 tcjswg = 0
+ tvoff = 0 tvfbsdoff = 0 saref = 3E-6
+ sbref = 3E-6 wlod = 0 ku0 = 7E-8
+ kvsat = 0.4 kvth0 = 3.5E-8 tku0 = 0
+ llodku0 = 0 wlodku0 = 1 llodvth = 0
+ wlodvth = 1 lku0 = 0 wku0 = 0
+ pku0 = 0 lkvth0 = 0 wkvth0 = 6.5E-7
+ pkvth0 = 0 stk2 = 0 lodk2 = 1
+ steta0 = 0 lodeta0 = 1

.model phv_model.31 pmos
+ level = 54 lmin = 2E-6 lmax = 4E-6 wmin = 1E-6
+ wmax = 3E-6 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 1.175E-8
+ toxm = 1.175E-8 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 1E23 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {1.2277E-8+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {4.5375E-8-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = -4.7338E-9 dwb = 0 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = -0.979159 lvth0 = -8.514514E-8
+ wvth0 = 2.290555E-8 pvth0 = 1.193942E-13 k1 = 0.595962
+ lk1 = -7.501062E-8 wk1 = 1.973425E-8 pk1 = 3.086927E-14
+ k2 = 3.12886E-2 lk2 = -5.322168E-9 wk2 = -1.761465E-8
+ pk2 = 2.670439E-14 k3 = -2.2405 k3b = -0.172
+ w0 = 0 lpe0 = 0 lpeb = 0
+ vbm = -3 dvtp0 = 0 dvtp1 = 0
+ dvt0 = 4.657 dvt1 = 0.34864 dvt2 = -0.030206
+ dvt0w = -2.2 dvt1w = 1.0163E6 dvt2w = 0
+ vfbsdoff = 0 u0 = 2.03004E-2 lu0 = 6.318867E-9
+ wu0 = -1.547121E-9 pu0 = -9.465007E-15 ua = 3.824629E-9
+ lua = -1.461103E-15 wua = -1.518719E-15 pua = 2.775247E-22
+ ub = -2.547604E-18 lub = 5.944632E-24 wub = 2.667101E-24
+ pub = -5.066726E-30 uc = -5.893907E-11 luc = 1.239993E-16
+ wuc = 1.194959E-17 puc = -5.694284E-23 ud = 0
+ up = 0 lp = 1 eu = 1.67
+ vsat = 6.497406E4 lvsat = 0.243228 wvsat = 0.146239
+ pvsat = -5.982357E-7 a0 = 0.846188 la0 = 1.445262E-7
+ wa0 = -5.283112E-8 pa0 = 1.468413E-13 ags = 0.35953
+ lags = -7.959178E-7 wags = -7.377186E-7 pags = 2.815343E-12
+ b0 = 0 b1 = 0 keta = -5.16874E-2
+ lketa = 1.570304E-7 wketa = 1.38656E-7 pketa = -5.355916E-13
+ a1 = 0 a2 = 0.5 rdsw = 788.47
+ rdswmin = 0 rdw = 0 rdwmin = 0
+ rsw = 0 rswmin = 0 prwb = 0.053538
+ prwg = 0 wr = 1 voff = -4.29193E-2
+ lvoff = -1.798537E-7 wvoff = -6.298346E-8 pvoff = 2.151629E-13
+ voffl = 0 minv = 0 nfactor = 2.623552
+ lnfactor = -3.26753E-6 wnfactor = -9.602857E-7 pnfactor = 3.26702E-12
+ eta0 = -4.78573E-2 leta0 = 4.998261E-7 weta0 = 1.992127E-7
+ peta0 = -7.787722E-13 etab = -0.115669 letab = 1.785308E-7
+ wetab = -2.00321E-8 petab = 7.831047E-14 dsub = 0.799307
+ ldsub = -9.35512E-7 wdsub = 4.59242E-8 pdsub = -1.795292E-13
+ cit = 8.578071E-6 lcit = 5.558677E-12 wcit = 4.230874E-12
+ pcit = -1.653954E-17 cdsc = 0 cdscb = 0
+ cdscd = 0 pclm = 1.575575 lpclm = -3.060287E-6
+ wpclm = -1.567491E-6 ppclm = 6.588659E-12 pdiblc1 = 0.675414
+ lpdiblc1 = -1.115756E-6 wpdiblc1 = -2.79252E-7 ppdiblc1 = 1.091666E-12
+ pdiblc2 = -2.315262E-3 lpdiblc2 = 1.409387E-8 wpdiblc2 = 3.516738E-9
+ ppdiblc2 = -1.374781E-14 pdiblcb = 0.259044 lpdiblcb = -1.110397E-6
+ wpdiblcb = -2.770691E-7 ppdiblcb = 1.083132E-12 drout = -2.85794E-2
+ ldrout = 2.300904E-6 wdrout = 5.014949E-7 pdrout = -1.960469E-12
+ pscbe1 = -3.026019E8 lpscbe1 = 1.335431E3 wpscbe1 = 435.699068
+ ppscbe1 = -9.93789E-4 pscbe2 = 1.057471E-7 lpscbe2 = -1.743405E-13
+ wpscbe2 = -8.828871E-14 ppscbe2 = 1.69188E-19 pvag = 0
+ delta = 0.01 fprout = 0 pdits = 0
+ pditsl = 0 pditsd = 0 lambda = 0
+ vtl = 0 lc = 5E-9 xn = 3
+ alpha0 = 2.14435E-4 lalpha0 = -7.071725E-10 walpha0 = -5.069323E-10
+ palpha0 = 1.853837E-15 alpha1 = -2.373533E-10 lalpha1 = 7.372103E-16
+ walpha1 = 4.221885E-16 palpha1 = -1.083132E-21 beta0 = 127.321069
+ lbeta0 = -2.861015E-4 wbeta0 = -1.7001E-4 pbeta0 = 4.696194E-10
+ aigbacc = 0.43 bigbacc = 0.054 cigbacc = 0.075
+ nigbacc = 1 aigbinv = 0.35 bigbinv = 0.03
+ cigbinv = 6E-3 eigbinv = 1.1 nigbinv = 3
+ aigc = 0.43 bigc = 0.054 cigc = 0.075
+ aigsd = 0.43 bigsd = 0.054 cigsd = 0.075
+ dlcig = 0 nigc = 1 poxedge = 1
+ pigcd = 1 ntox = 1 toxref = 1.175E-8
+ agidl = 6.988925E-10 lagidl = -1.212567E-14 wagidl = 2.613367E-14
+ pagidl = 3.512544E-20 bgidl = 3.025185E9 lbgidl = -3.805331E3
+ wbgidl = -1.638883E3 pbgidl = 4.197138E-3 cgidl = 1.175864E3
+ lcgidl = -1.696329E-3 wcgidl = -9.911252E-4 pcgidl = 2.921479E-9
+ egidl = -3.586751 legidl = 1.117207E-5 wegidl = 5.955142E-6
+ pegidl = -1.287414E-11 noia = 3E40 noib = 8.53E24
+ noic = 8.4E7 em = 4.1E7 af = 1
+ ef = 0.88 kf = 0 lintnoi = 0
+ tnoia = 1.5 tnoib = 3.5 ntnoi = 1
+ rnoia = 0.577 rnoib = 0.37 xpart = 0
+ cgso = {1.94171E-10/sw_func_tox_hv_ratio} cgdo = {1.94171E-10/sw_func_tox_hv_ratio} cgbo = {0/sw_func_tox_hv_ratio}
+ ckappas = 0.6 cf = 1.2E-11 clc = 1E-7
+ cle = 0.6 dlc = 4.4983E-8 dwc = 0
+ vfbcv = -0.144689 noff = 4 voffcv = 0
+ acde = 0.401 moin = 15.773 cgsl = {9.82591E-12/sw_func_tox_hv_ratio}
+ cgdl = {9.82591E-12/sw_func_tox_hv_ratio} ijthsrev = 0.1 ijthsfwd = 0.1
+ xjbvs = 1 bvs = 12.69 jss = 2.1483E-5
+ jsws = 4.02E-12 cjs = {sw_psd_nw_cj} mjs = 0.33956
+ mjsws = 0.24676 cjsws = {9.960545E-11*sw_func_psd_nw_cj} cjswgs = {1.47314E-10*sw_func_psd_nw_cj}
+ mjswgs = 0.81 pbs = 0.6587 pbsws = 1
+ pbswgs = 3 xrcrg1 = 12 xrcrg2 = 1
+ rbpb = 50 rbpd = 50 rbps = 50
+ rbdb = 50 rbsb = 50 gbmin = 1E-12
+ tnom = 30 ute = -1.775057 lute = 5.781633E-7
+ wute = 3.495578E-7 pute = -5.399415E-13 kt1 = -0.595578
+ lkt1 = 7.653658E-8 wkt1 = 5.541382E-8 pkt1 = -2.166265E-13
+ kt1l = 0 kt2 = -0.019032 ua1 = -3.812681E-10
+ lua1 = 1.576851E-15 wua1 = -3.06106E-16 pua1 = 1.196645E-21
+ ub1 = -4.077704E-18 lub1 = -1.314192E-24 wub1 = 2.010204E-24
+ pub1 = -1.781753E-31 uc1 = -1.092E-10 at = 2.223866E5
+ lat = 4.75188E-2 wat = 0.186188 pat = -7.846428E-7
+ prt = 0 njs = 1.3632 xtis = 10
+ tpb = 1.671E-3 tpbsw = 0 tpbswg = 0
+ tcj = 9.6E-4 tcjsw = 3E-5 tcjswg = 0
+ tvoff = 0 tvfbsdoff = 0 saref = 3E-6
+ sbref = 3E-6 wlod = 0 ku0 = 7E-8
+ kvsat = 0.4 kvth0 = 3.5E-8 tku0 = 0
+ llodku0 = 0 wlodku0 = 1 llodvth = 0
+ wlodvth = 1 lku0 = 0 wku0 = 0
+ pku0 = 0 lkvth0 = 0 wkvth0 = 6.5E-7
+ pkvth0 = 0 stk2 = 0 lodk2 = 1
+ steta0 = 0 lodeta0 = 1

.model phv_model.32 pmos
+ level = 54 lmin = 1E-6 lmax = 2E-6 wmin = 1E-6
+ wmax = 3E-6 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 1.175E-8
+ toxm = 1.175E-8 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 1E23 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {1.2277E-8+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {4.5375E-8-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = -4.7338E-9 dwb = 0 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = -1.06634 lvth0 = 8.13056E-8
+ wvth0 = 1.106423E-7 pvth0 = -4.811719E-14 k1 = 0.543505
+ lk1 = 2.514315E-8 wk1 = 4.627378E-8 pk1 = -1.980131E-14
+ k2 = 2.20795E-2 lk2 = 1.226043E-8 wk2 = 2.548511E-9
+ pk2 = -1.179213E-14 k3 = -2.2405 k3b = -0.172
+ w0 = 0 lpe0 = 0 lpeb = 0
+ vbm = -3 dvtp0 = 0 dvtp1 = 0
+ dvt0 = 4.657 dvt1 = 0.34864 dvt2 = -0.030206
+ dvt0w = -2.2 dvt1w = 1.0163E6 dvt2w = 0
+ vfbsdoff = 0 u0 = 2.85264E-2 lu0 = -9.386587E-9
+ wu0 = -9.58644E-9 pu0 = 5.884063E-15 ua = 4.025692E-9
+ lua = -1.844984E-15 wua = -1.680917E-15 pua = 5.872014E-22
+ ub = 7.745995E-19 lub = -3.982854E-25 wub = -7.690582E-25
+ pub = 1.493762E-30 uc = 1.127653E-11 luc = -1.005981E-17
+ wuc = -3.196879E-17 puc = 2.690832E-23 ud = 0
+ up = 0 lp = 1 eu = 1.67
+ vsat = 3.22856E5 lvsat = -0.249133 wvsat = -0.316409
+ pvsat = 2.850759E-7 a0 = 1.002577 la0 = -1.540602E-7
+ wa0 = 1.021598E-8 pa0 = 2.646866E-14 ags = -0.74749
+ lags = 1.317659E-6 wags = 1.404499E-6 pags = -1.274686E-12
+ b0 = 0 b1 = 0 keta = 0.134109
+ lketa = -1.977022E-7 wketa = -2.672183E-7 pketa = 2.393238E-13
+ a1 = 0 a2 = 0.5 rdsw = 788.47
+ rdswmin = 0 rdw = 0 rdwmin = 0
+ rsw = 0 rswmin = 0 prwb = 0.053538
+ prwg = 0 wr = 1 voff = -0.191935
+ lvoff = 1.046555E-7 wvoff = 9.74041E-8 pvoff = -9.105704E-14
+ voffl = 0 minv = 0 nfactor = 0.19865
+ lnfactor = 1.362213E-6 wnfactor = 1.493473E-6 pnfactor = -1.417819E-12
+ eta0 = 0.41412 leta0 = -3.822041E-7 weta0 = -4.390225E-7
+ peta0 = 4.397783E-13 etab = -4.26585E-2 letab = 3.913589E-8
+ wetab = 4.110153E-8 petab = -3.84089E-14 dsub = 0.322667
+ ldsub = -2.548601E-8 wdsub = -1.036237E-7 pdsub = 1.059952E-13
+ cit = 1.739011E-5 lcit = -1.126571E-11 wcit = -8.461747E-12
+ pcit = 7.693844E-18 cdsc = 0 cdscb = 0
+ cdscd = 0 pclm = -1.1173 lpclm = 2.081085E-6
+ wpclm = 3.510382E-6 ppclm = -3.10627E-12 pdiblc1 = -0.22243
+ lpdiblc1 = 5.984528E-7 wpdiblc1 = 6.565129E-7 ppdiblc1 = -6.949433E-13
+ pdiblc2 = 8.528579E-3 lpdiblc2 = -6.609733E-9 wpdiblc2 = -7.701825E-9
+ ppdiblc2 = 7.671232E-15 pdiblcb = -0.593087 lpdiblcb = 5.165331E-7
+ wpdiblcb = 5.541382E-7 ppdiblcb = -5.038502E-13 drout = 2.134256
+ ldrout = -1.82849E-6 wdrout = -1.780583E-6 pdrout = 2.396589E-12
+ pscbe1 = 4.905104E8 lpscbe1 = -178.819075 wpscbe1 = -177.179467
+ ppscbe1 = 1.763494E-4 pscbe2 = 1.426307E-8 lpscbe2 = 3.254309E-16
+ wpscbe2 = 8.024358E-16 ppscbe2 = -9.092934E-22 pvag = 0
+ delta = 0.01 fprout = 0 pdits = 0
+ pditsl = 0 pditsd = 0 lambda = 0
+ vtl = 0 lc = 5E-9 xn = 3
+ alpha0 = -3.565746E-4 lalpha0 = 3.830277E-10 walpha0 = 8.775056E-10
+ palpha0 = -7.894012E-16 alpha1 = 2.840435E-10 lalpha1 = -2.582666E-16
+ walpha1 = -2.770691E-16 palpha1 = 2.519251E-22 beta0 = -88.704544
+ lbeta0 = 1.263454E-4 wbeta0 = 1.452933E-4 pbeta0 = -1.323734E-10
+ aigbacc = 0.43 bigbacc = 0.054 cigbacc = 0.075
+ nigbacc = 1 aigbinv = 0.35 bigbinv = 0.03
+ cigbinv = 6E-3 eigbinv = 1.1 nigbinv = 3
+ aigc = 0.43 bigc = 0.054 cigc = 0.075
+ aigsd = 0.43 bigsd = 0.054 cigsd = 0.075
+ dlcig = 0 nigc = 1 poxedge = 1
+ pigcd = 1 ntox = 1 toxref = 1.175E-8
+ agidl = -1.809264E-8 lagidl = 2.375207E-14 wagidl = 9.047437E-14
+ pagidl = -8.771704E-20 bgidl = 5.393949E8 lbgidl = 940.664357
+ wbgidl = 1.095547E3 pbgidl = -1.023572E-3 cgidl = -536.078606
+ lcgidl = 1.572198E-3 wcgidl = 1.767854E-3 pcgidl = -2.346103E-9
+ egidl = 3.31468 legidl = -2.004484E-6 wegidl = -6.083788E-7
+ pegidl = -3.42743E-13 noia = 3E40 noib = 8.53E24
+ noic = 8.4E7 em = 4.1E7 af = 1
+ ef = 0.88 kf = 0 lintnoi = 0
+ tnoia = 1.5 tnoib = 3.5 ntnoi = 1
+ rnoia = 0.577 rnoib = 0.37 xpart = 0
+ cgso = {1.94171E-10/sw_func_tox_hv_ratio} cgdo = {1.94171E-10/sw_func_tox_hv_ratio} cgbo = {0/sw_func_tox_hv_ratio}
+ ckappas = 0.6 cf = 1.2E-11 clc = 1E-7
+ cle = 0.6 dlc = 4.4983E-8 dwc = 0
+ vfbcv = -0.144689 noff = 4 voffcv = 0
+ acde = 0.401 moin = 15.773 cgsl = {9.82591E-12/sw_func_tox_hv_ratio}
+ cgdl = {9.82591E-12/sw_func_tox_hv_ratio} ijthsrev = 0.1 ijthsfwd = 0.1
+ xjbvs = 1 bvs = 12.69 jss = 2.1483E-5
+ jsws = 4.02E-12 cjs = {sw_psd_nw_cj} mjs = 0.33956
+ mjsws = 0.24676 cjsws = {9.960545E-11*sw_func_psd_nw_cj} cjswgs = {1.47314E-10*sw_func_psd_nw_cj}
+ mjswgs = 0.81 pbs = 0.6587 pbsws = 1
+ pbswgs = 3 xrcrg1 = 12 xrcrg2 = 1
+ rbpb = 50 rbpd = 50 rbps = 50
+ rbdb = 50 rbsb = 50 gbmin = 1E-12
+ tnom = 30 ute = -1.477755 lute = 1.053796E-8
+ wute = 1.129373E-7 pute = -8.817378E-14 kt1 = -0.491292
+ lkt1 = -1.22573E-7 wkt1 = -1.002717E-7 pkt1 = 8.061603E-14
+ kt1l = 0 kt2 = -0.019032 ua1 = 3.466453E-10
+ lua1 = 1.870824E-16 wua1 = 6.122119E-16 pua1 = -5.566537E-22
+ ub1 = -5.834523E-18 lub1 = 2.040014E-24 wub1 = 3.659806E-24
+ pub1 = -3.327678E-30 uc1 = -1.092E-10 at = 4.44833E5
+ lat = -0.377187 wat = -0.429163 pat = 3.902168E-7
+ prt = 0 njs = 1.3632 xtis = 10
+ tpb = 1.671E-3 tpbsw = 0 tpbswg = 0
+ tcj = 9.6E-4 tcjsw = 3E-5 tcjswg = 0
+ tvoff = 0 tvfbsdoff = 0 saref = 3E-6
+ sbref = 3E-6 wlod = 0 ku0 = 7E-8
+ kvsat = 0.4 kvth0 = 3.5E-8 tku0 = 0
+ llodku0 = 0 wlodku0 = 1 llodvth = 0
+ wlodvth = 1 lku0 = 0 wku0 = 0
+ pku0 = 0 lkvth0 = 0 wkvth0 = 6.5E-7
+ pkvth0 = 0 stk2 = 0 lodk2 = 1
+ steta0 = 0 lodeta0 = 1

.model phv_model.33 pmos
+ level = 54 lmin = 8E-7 lmax = 1E-6 wmin = 1E-6
+ wmax = 3E-6 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 1.175E-8
+ toxm = 1.175E-8 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 1E23 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {1.2277E-8+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {4.5375E-8-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = -4.7338E-9 dwb = 0 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = -0.982717 lvth0 = 5.271448E-9
+ wvth0 = 7.497305E-8 pvth0 = -1.568491E-14 k1 = 0.537759
+ lk1 = 3.036744E-8 wk1 = 1.238711E-7 pk1 = -9.035668E-14
+ k2 = 4.92495E-2 lk2 = -1.244396E-8 wk2 = -5.114239E-8
+ pk2 = 3.702632E-14 k3 = -2.2405 k3b = -0.172
+ w0 = 0 lpe0 = 0 lpeb = 0
+ vbm = -3 dvtp0 = 0 dvtp1 = 0
+ dvt0 = 4.657 dvt1 = 0.34864 dvt2 = -0.030206
+ dvt0w = -2.2 dvt1w = 1.0163E6 dvt2w = 0
+ vfbsdoff = 0 u0 = 1.96893E-2 lu0 = -1.351485E-9
+ wu0 = -7.537726E-9 pu0 = 4.02127E-15 ua = 2.768587E-9
+ lua = -7.019615E-16 wua = -3.33222E-15 pua = 2.088648E-21
+ ub = -3.611362E-19 lub = 6.343822E-25 wub = 2.949756E-24
+ pub = -1.88757E-30 uc = 7.86919E-13 luc = -5.221297E-19
+ wuc = -4.08344E-18 puc = 1.553569E-24 ud = 0
+ up = 0 lp = 1 eu = 1.67
+ vsat = 6.777173E4 lvsat = -1.71981E-2 wvsat = -0.05916
+ pvsat = 5.117201E-8 a0 = 0.699189 la0 = 1.217949E-7
+ wa0 = 4.378903E-7 pa0 = -3.623942E-13 ags = 0.75599
+ lags = -4.937942E-8 wags = -1.590001E-7 pags = 1.469258E-13
+ b0 = 0 b1 = 0 keta = -4.38609E-2
+ lketa = -3.588264E-8 wketa = -1.214312E-7 pketa = 1.067669E-13
+ a1 = 0 a2 = 0.5 rdsw = 788.47
+ rdswmin = 0 rdw = 0 rdwmin = 0
+ rsw = 0 rswmin = 0 prwb = 0.053538
+ prwg = 0 wr = 1 voff = -8.37017E-2
+ lvoff = 6.244003E-9 wvoff = 1.769187E-8 pvoff = -1.857869E-14
+ voffl = 0 minv = 0 nfactor = 1.607474
+ lnfactor = 8.124037E-8 wnfactor = 1.999973E-7 pnfactor = -2.417263E-13
+ eta0 = -6.28192E-2 leta0 = 5.145292E-8 weta0 = 2.130245E-7
+ peta0 = -1.530954E-13 etab = -5.338636E-3 letab = 5.202787E-9
+ wetab = 1.588482E-8 petab = -1.548061E-14 dsub = 0.22077
+ ldsub = 6.716342E-8 wdsub = 2.327374E-7 pdsub = -1.998411E-13
+ cit = 1.364794E-5 lcit = -7.863138E-12 wcit = -2.573147E-11
+ pcit = 2.339634E-17 cdsc = 0 cdscb = 0
+ cdscd = 0 pclm = 0.972135 lpclm = 1.812658E-7
+ wpclm = 6.872604E-7 ppclm = -5.393465E-13 pdiblc1 = 0.658671
+ lpdiblc1 = -2.026881E-7 wpdiblc1 = -7.710712E-7 ppdiblc1 = 6.030876E-13
+ pdiblc2 = 9.199472E-3 lpdiblc2 = -7.219743E-9 wpdiblc2 = -2.289096E-8
+ ppdiblc2 = 2.148195E-14 pdiblcb = -0.025 drout = -0.661793
+ ldrout = 7.138177E-7 wdrout = 3.191113E-6 pdrout = -2.123926E-12
+ pscbe1 = 3.939577E8 lpscbe1 = -91.028451 wpscbe1 = -281.112258
+ ppscbe1 = 2.708502E-4 pscbe2 = 1.300548E-8 lpscbe2 = 1.468894E-15
+ wpscbe2 = 4.609223E-15 ppscbe2 = -4.370615E-21 pvag = 0
+ delta = 0.01 fprout = 0 pdits = 0
+ pditsl = 0 pditsd = 0 lambda = 0
+ vtl = 0 lc = 5E-9 xn = 3
+ alpha0 = -7.57516E-6 lalpha0 = 6.569994E-11 walpha0 = 2.243139E-10
+ palpha0 = -1.954866E-16 alpha1 = 0 beta0 = 45.919938
+ lbeta0 = 3.938064E-6 wbeta0 = 1.259502E-5 pbeta0 = -1.17175E-11
+ aigbacc = 0.43 bigbacc = 0.054 cigbacc = 0.075
+ nigbacc = 1 aigbinv = 0.35 bigbinv = 0.03
+ cigbinv = 6E-3 eigbinv = 1.1 nigbinv = 3
+ aigc = 0.43 bigc = 0.054 cigc = 0.075
+ aigsd = 0.43 bigsd = 0.054 cigsd = 0.075
+ dlcig = 0 nigc = 1 poxedge = 1
+ pigcd = 1 ntox = 1 toxref = 1.175E-8
+ agidl = 1.818897E-8 lagidl = -9.236986E-15 wagidl = -3.622477E-14
+ pagidl = 2.748415E-20 bgidl = 1.998731E9 lbgidl = -386.23734
+ wbgidl = -1.294115E3 pbgidl = 1.149228E-3 cgidl = 1.452164E3
+ lcgidl = -2.356111E-4 wcgidl = -1.583425E-3 pcgidl = 7.01048E-10
+ egidl = 1.217569 legidl = -9.768645E-8 wegidl = -1.305001E-6
+ pegidl = 2.906608E-13 noia = 3E40 noib = 8.53E24
+ noic = 8.4E7 em = 4.1E7 af = 1
+ ef = 0.88 kf = 0 lintnoi = 0
+ tnoia = 1.5 tnoib = 3.5 ntnoi = 1
+ rnoia = 0.577 rnoib = 0.37 xpart = 0
+ cgso = {1.94171E-10/sw_func_tox_hv_ratio} cgdo = {1.94171E-10/sw_func_tox_hv_ratio} cgbo = {0/sw_func_tox_hv_ratio}
+ ckappas = 0.6 cf = 1.2E-11 clc = 1E-7
+ cle = 0.6 dlc = 4.4983E-8 dwc = 0
+ vfbcv = -0.144689 noff = 4 voffcv = 0
+ acde = 0.401 moin = 15.773 cgsl = {9.82591E-12/sw_func_tox_hv_ratio}
+ cgdl = {9.82591E-12/sw_func_tox_hv_ratio} ijthsrev = 0.1 ijthsfwd = 0.1
+ xjbvs = 1 bvs = 12.69 jss = 2.1483E-5
+ jsws = 4.02E-12 cjs = {sw_psd_nw_cj} mjs = 0.33956
+ mjsws = 0.24676 cjsws = {9.960545E-11*sw_func_psd_nw_cj} cjswgs = {1.47314E-10*sw_func_psd_nw_cj}
+ mjswgs = 0.81 pbs = 0.6587 pbsws = 1
+ pbswgs = 3 xrcrg1 = 12 xrcrg2 = 1
+ rbpb = 50 rbpd = 50 rbps = 50
+ rbdb = 50 rbsb = 50 gbmin = 1E-12
+ tnom = 30 ute = -1.518053 lute = 4.717883E-8
+ wute = 1.70352E-7 pute = -1.403781E-13 kt1 = -0.630422
+ lkt1 = 3.931569E-9 wkt1 = 1.256189E-9 pkt1 = -1.169817E-14
+ kt1l = 0 kt2 = -0.019032 ua1 = 5.524E-10
+ ub1 = -3.5909E-18 uc1 = -1.092E-10 at = 1.270412E4
+ lat = 1.57263E-2 wat = 5.14629E-2 pat = -4.679269E-8
+ prt = 0 njs = 1.3632 xtis = 10
+ tpb = 1.671E-3 tpbsw = 0 tpbswg = 0
+ tcj = 9.6E-4 tcjsw = 3E-5 tcjswg = 0
+ tvoff = 0 tvfbsdoff = 0 saref = 2.81E-6
+ sbref = 2.81E-6 wlod = 0 ku0 = 7E-8
+ kvsat = 0.4 kvth0 = 3.5E-8 tku0 = 0
+ llodku0 = 0 wlodku0 = 1 llodvth = 0
+ wlodvth = 1 lku0 = 0 wku0 = 0
+ pku0 = 0 lkvth0 = 0 wkvth0 = 6.5E-7
+ pkvth0 = 0 stk2 = 0 lodk2 = 1
+ steta0 = 0 lodeta0 = 1

.model phv_model.34 pmos
+ level = 54 lmin = 6E-7 lmax = 8E-7 wmin = 1E-6
+ wmax = 3E-6 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 1.175E-8
+ toxm = 1.175E-8 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 1E23 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {1.2277E-8+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {4.5375E-8-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = -4.7338E-9 dwb = 0 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = -1.008005 lvth0 = 2.320703E-8
+ wvth0 = 7.221912E-8 pvth0 = -1.373168E-14 k1 = 0.654744
+ lk1 = -5.26045E-8 wk1 = -2.010296E-7 pk1 = 1.400791E-13
+ k2 = -9.686102E-3 lk2 = 2.935614E-8 wk2 = 6.27013E-8
+ pk2 = -4.371731E-14 k3 = -2.2405 k3b = -0.172
+ w0 = 0 lpe0 = 0 lpeb = 0
+ vbm = -3 dvtp0 = 0 dvtp1 = 0
+ dvt0 = 4.657 dvt1 = 0.34864 dvt2 = -0.030206
+ dvt0w = -2.2 dvt1w = 1.0163E6 dvt2w = 0
+ vfbsdoff = 0 u0 = 1.49618E-2 lu0 = 2.001509E-9
+ wu0 = 3.549781E-9 pu0 = -3.842545E-15 ua = -1.081638E-9
+ lua = 2.028811E-15 wua = 2.851975E-15 pua = -2.297492E-21
+ ub = 4.232191E-18 lub = -2.623435E-24 wub = -3.362438E-24
+ pub = 2.589354E-30 uc = 6.100663E-12 luc = -4.290903E-18
+ wuc = -5.648311E-18 puc = 2.663454E-24 ud = 0
+ up = 0 lp = 1 eu = 1.67
+ vsat = -3.590138E4 lvsat = 0.056332 wvsat = 5.39342E-2
+ pvsat = -2.904001E-8 a0 = 0.938825 la0 = -4.816662E-8
+ wa0 = -2.535599E-7 pa0 = 1.280169E-13 ags = 0.599221
+ lags = 6.180833E-8 wags = 1.6678E-7 pags = -8.413377E-14
+ b0 = 0 b1 = 0 keta = -0.235907
+ lketa = 1.003264E-7 wketa = 1.344658E-7 pketa = -7.472808E-14
+ a1 = 0 a2 = 0.5 rdsw = 788.47
+ rdswmin = 0 rdw = 0 rdwmin = 0
+ rsw = 0 rswmin = 0 prwb = 0.053538
+ prwg = 0 wr = 1 voff = -8.90607E-2
+ lvoff = 1.004488E-8 wvoff = -3.747237E-9 pvoff = -3.373008E-15
+ voffl = 0 minv = 0 nfactor = 1.518852
+ lnfactor = 1.440953E-7 wnfactor = -2.15977E-7 pnfactor = 5.330345E-14
+ eta0 = 5.57775E-2 leta0 = -3.266181E-8 weta0 = -7.520594E-8
+ peta0 = 5.133204E-14 etab = 7.081797E-3 letab = -3.606405E-9
+ wetab = -2.10715E-8 petab = 1.073066E-14 dsub = 0.415237
+ ldsub = -7.076193E-8 wdsub = -1.627735E-7 pdsub = 8.067493E-14
+ cit = -1.637919E-5 lcit = 1.34336E-11 wcit = 2.573147E-11
+ pcit = -1.310375E-17 cdsc = 0 cdscb = 0
+ cdscd = 0 pclm = 2.036813 lpclm = -5.73857E-7
+ wpclm = -7.312609E-7 ppclm = 4.667397E-13 pdiblc1 = 8.63172E-2
+ lpdiblc1 = 2.032539E-7 wpdiblc1 = 4.968274E-7 ppdiblc1 = -2.961695E-13
+ pdiblc2 = -3.69548E-2 lpdiblc2 = 2.551519E-8 wpdiblc2 = 3.939806E-8
+ ppdiblc2 = -2.269653E-14 pdiblcb = -0.025 drout = 0.384149
+ ldrout = -2.80162E-8 wdrout = -8.093243E-8 pdrout = 1.967722E-13
+ pscbe1 = -1.529191E8 lpscbe1 = 296.843914 wpscbe1 = 584.529801
+ ppscbe1 = -3.431064E-4 pscbe2 = 2.046211E-8 lpscbe2 = -3.81972E-15
+ wpscbe2 = -9.615305E-15 ppscbe2 = 5.718132E-21 pvag = 0
+ delta = 0.01 fprout = 0 pdits = 0
+ pditsl = 0 pditsd = 0 lambda = 0
+ vtl = 0 lc = 5E-9 xn = 3
+ alpha0 = 2.731563E-4 lalpha0 = -1.334088E-10 walpha0 = -2.278348E-10
+ palpha0 = 1.251999E-16 alpha1 = 0 beta0 = 70.582212
+ lbeta0 = -1.355365E-5 wbeta0 = -2.43734E-5 pbeta0 = 1.450236E-11
+ aigbacc = 0.43 bigbacc = 0.054 cigbacc = 0.075
+ nigbacc = 1 aigbinv = 0.35 bigbinv = 0.03
+ cigbinv = 6E-3 eigbinv = 1.1 nigbinv = 3
+ aigc = 0.43 bigc = 0.054 cigc = 0.075
+ aigsd = 0.43 bigsd = 0.054 cigsd = 0.075
+ dlcig = 0 nigc = 1 poxedge = 1
+ pigcd = 1 ntox = 1 toxref = 1.175E-8
+ agidl = 3.238713E-8 lagidl = -1.930703E-14 wagidl = -1.215006E-13
+ pagidl = 8.796602E-20 bgidl = 2.339548E8 lbgidl = 865.430452
+ wbgidl = 2.112071E3 pbgidl = -1.266609E-3 cgidl = 3.201503E3
+ lcgidl = -1.47633E-3 wcgidl = -3.757996E-3 pcgidl = 2.243363E-9
+ egidl = 3.513778 legidl = -1.726273E-6 wegidl = -5.879968E-6
+ pegidl = 3.535456E-12 noia = 3E40 noib = 8.53E24
+ noic = 8.4E7 em = 4.1E7 af = 1
+ ef = 0.88 kf = 0 lintnoi = 0
+ tnoia = 1.5 tnoib = 3.5 ntnoi = 1
+ rnoia = 0.577 rnoib = 0.37 xpart = 0
+ cgso = {1.94171E-10/sw_func_tox_hv_ratio} cgdo = {1.94171E-10/sw_func_tox_hv_ratio} cgbo = {0/sw_func_tox_hv_ratio}
+ ckappas = 0.6 cf = 1.2E-11 clc = 1E-7
+ cle = 0.6 dlc = 4.4983E-8 dwc = 0
+ vfbcv = -0.144689 noff = 4 voffcv = 0
+ acde = 0.401 moin = 15.773 cgsl = {9.82591E-12/sw_func_tox_hv_ratio}
+ cgdl = {9.82591E-12/sw_func_tox_hv_ratio} ijthsrev = 0.1 ijthsfwd = 0.1
+ xjbvs = 1 bvs = 12.69 jss = 2.1483E-5
+ jsws = 4.02E-12 cjs = {sw_psd_nw_cj} mjs = 0.33956
+ mjsws = 0.24676 cjsws = {9.960545E-11*sw_func_psd_nw_cj} cjswgs = {1.47314E-10*sw_func_psd_nw_cj}
+ mjswgs = 0.81 pbs = 0.6587 pbsws = 1
+ pbswgs = 3 xrcrg1 = 12 xrcrg2 = 1
+ rbpb = 50 rbpd = 50 rbps = 50
+ rbdb = 50 rbsb = 50 gbmin = 1E-12
+ tnom = 30 ute = -1.292669 lute = -1.126743E-7
+ wute = -5.267809E-7 pute = 3.540634E-13 kt1 = -0.582358
+ lkt1 = -3.015774E-8 wkt1 = -2.447528E-8 pkt1 = 6.551877E-15
+ kt1l = 0 kt2 = -0.019032 ua1 = 5.524E-10
+ ub1 = -2.558271E-18 lub1 = -7.323919E-25 wub1 = -5.282517E-24
+ pub1 = 3.746625E-30 uc1 = -3.656705E-10 luc1 = 1.819017E-16
+ wuc1 = 2.501731E-16 puc1 = -1.774353E-22 at = 6.791596E4
+ lat = -2.34327E-2 wat = -2.19021E-2 pat = 5.241501E-9
+ prt = 0 njs = 1.3632 xtis = 10
+ tpb = 1.671E-3 tpbsw = 0 tpbswg = 0
+ tcj = 9.6E-4 tcjsw = 3E-5 tcjswg = 0
+ tvoff = 0 tvfbsdoff = 0 saref = 2.41E-6
+ sbref = 2.41E-6 wlod = 0 ku0 = 7E-8
+ kvsat = 0.4 kvth0 = 3.5E-8 tku0 = 0
+ llodku0 = 0 wlodku0 = 1 llodvth = 0
+ wlodvth = 1 lku0 = 0 wku0 = 0
+ pku0 = 0 lkvth0 = 0 wkvth0 = 6.5E-7
+ pkvth0 = 0 stk2 = 0 lodk2 = 1
+ steta0 = 0 lodeta0 = 1

.model phv_model.35 pmos
+ level = 54 lmin = 5E-7 lmax = 6E-7 wmin = 1E-6
+ wmax = 3E-6 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 1.175E-8
+ toxm = 1.175E-8 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 1E23 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {1.2277E-8+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {4.5375E-8-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = -4.7338E-9 dwb = 0 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = -0.730216 lvth0 = -1.182573E-7
+ wvth0 = -5.358002E-8 pvth0 = 5.033153E-14 k1 = 0.462169
+ lk1 = 4.546439E-8 wk1 = 4.321028E-7 pk1 = -1.823435E-13
+ k2 = 7.56535E-2 lk2 = -1.410308E-8 wk2 = -1.40105E-7
+ pk2 = 5.95618E-14 k3 = -2.2405 k3b = -0.172
+ w0 = 0 lpe0 = 0 lpeb = 0
+ vbm = -3 dvtp0 = 0 dvtp1 = 0
+ dvt0 = 4.657 dvt1 = 0.34864 dvt2 = -0.030206
+ dvt0w = -2.2 dvt1w = 1.0163E6 dvt2w = 0
+ vfbsdoff = 0 u0 = 6.04869E-3 lu0 = 6.540505E-9
+ wu0 = 5.089661E-9 pu0 = -4.626728E-15 ua = 1.486048E-9
+ lua = 7.212167E-16 wua = -6.06195E-16 pua = -5.36419E-22
+ ub = -3.940762E-18 lub = 1.538641E-24 wub = 3.539184E-24
+ pub = -9.252973E-31 uc = 1.954697E-10 luc = -1.007271E-16
+ wuc = -1.806001E-16 puc = 9.175763E-23 ud = 0
+ up = 0 lp = 1 eu = 1.67
+ vsat = -1.420898E5 lvsat = 0.110408 wvsat = 3.53244E-2
+ pvsat = -1.956299E-8 a0 = 0.101406 la0 = 3.782889E-7
+ wa0 = 1.20653E-6 pa0 = -6.155341E-13 ags = 2.743907
+ lags = -1.030373E-6 wags = 4.48761E-7 pags = -2.277326E-13
+ b0 = 0 b1 = 0 keta = -0.209552
+ lketa = 8.690489E-8 wketa = -1.745173E-8 pketa = 2.635921E-15
+ a1 = 0 a2 = 0.5 rdsw = 788.47
+ rdswmin = 0 rdw = 0 rdwmin = 0
+ rsw = 0 rswmin = 0 prwb = 0.053538
+ prwg = 0 wr = 1 voff = 0.154131
+ lvoff = -1.138004E-7 wvoff = -9.575661E-8 pvoff = 4.348277E-14
+ voffl = 0 minv = 0 nfactor = 2.593255
+ lnfactor = -4.030443E-7 wnfactor = -5.855958E-7 pnfactor = 2.415318E-13
+ eta0 = -0.605863 leta0 = 3.042787E-7 weta0 = 5.532445E-8
+ peta0 = -1.514056E-14 etab = 7.01369E-2 letab = -3.57172E-8
+ wetab = -2.471816E-8 petab = 1.258772E-14 dsub = 0.177416
+ ldsub = 5.034817E-8 wdsub = 6.661531E-8 pdsub = -3.614131E-14
+ cit = 1.996811E-8 lcit = 5.082331E-12 wcit = 2.969505E-11
+ pcit = -1.51222E-17 cdsc = 0 cdscb = 0
+ cdscd = 0 pclm = 2.22514 lpclm = -6.697625E-7
+ wpclm = 7.350933E-7 ppclm = -2.800012E-13 pdiblc1 = 1.584456
+ lpdiblc1 = -5.596733E-7 wpdiblc1 = -9.594231E-8 ppdiblc1 = 5.698469E-15
+ pdiblc2 = 4.77972E-2 lpdiblc2 = -1.764477E-8 wpdiblc2 = -1.59344E-8
+ ppdiblc2 = 5.481521E-15 pdiblcb = 0.7935 lpdiblcb = -4.168211E-7
+ drout = -2.416386 ldrout = 1.398156E-6 wdrout = 1.555574E-6
+ pdrout = -6.366186E-13 pscbe1 = 1.543823E9 lpscbe1 = -567.222029
+ wpscbe1 = -3.01794E3 ppscbe1 = 1.491451E-3 pscbe2 = -1.118928E-8
+ lpscbe2 = 1.229875E-14 wpscbe2 = 6.0814E-14 ppscbe2 = -3.014799E-20
+ pvag = 0 delta = 0.01 fprout = 0
+ pdits = 0 pditsl = 0 pditsd = 0
+ lambda = 0 vtl = 0 lc = 5E-9
+ xn = 3 alpha0 = 6.49439E-5 lalpha0 = -2.737668E-11
+ walpha0 = 6.799268E-11 palpha0 = -2.545031E-17 alpha1 = -6.088506E-10
+ lalpha1 = 3.100572E-16 walpha1 = 5.939009E-16 palpha1 = -3.02444E-22
+ beta0 = 281.663816 lbeta0 = -1.21047E-4 wbeta0 = -1.874921E-4
+ pbeta0 = 9.757054E-11 aigbacc = 0.43 bigbacc = 0.054
+ cigbacc = 0.075 nigbacc = 1 aigbinv = 0.35
+ bigbinv = 0.03 cigbinv = 6E-3 eigbinv = 1.1
+ nigbinv = 3 aigc = 0.43 bigc = 0.054
+ cigc = 0.075 aigsd = 0.43 bigsd = 0.054
+ cigsd = 0.075 dlcig = 0 nigc = 1
+ poxedge = 1 pigcd = 1 ntox = 1
+ toxref = 1.175E-8 agidl = -1.02631E-7 lagidl = 4.945097E-14
+ wagidl = 2.840806E-13 pagidl = -1.185762E-19 bgidl = 6.501561E9
+ lbgidl = -2.326348E3 wbgidl = -6.817177E3 pbgidl = 3.280611E-3
+ cgidl = -2.539371E3 lcgidl = 1.447211E-3 wcgidl = 6.077981E-3
+ pcgidl = -2.765609E-9 egidl = -11.275933 legidl = 5.805388E-6
+ wegidl = 1.64858E-5 pegidl = -7.85431E-12 noia = 3E40
+ noib = 8.53E24 noic = 8.4E7 em = 4.1E7
+ af = 1 ef = 0.88 kf = 0
+ lintnoi = 0 tnoia = 1.5 tnoib = 3.5
+ ntnoi = 1 rnoia = 0.577 rnoib = 0.37
+ xpart = 0 cgso = {1.94171E-10/sw_func_tox_hv_ratio} cgdo = {1.94171E-10/sw_func_tox_hv_ratio}
+ cgbo = {0/sw_func_tox_hv_ratio} ckappas = 0.6 cf = 1.2E-11
+ clc = 1E-7 cle = 0.6 dlc = 4.4983E-8
+ dwc = 0 vfbcv = -0.144689 noff = 4
+ voffcv = 0 acde = 0.401 moin = 15.773
+ cgsl = {9.82591E-12/sw_func_tox_hv_ratio} cgdl = {9.82591E-12/sw_func_tox_hv_ratio} ijthsrev = 0.1
+ ijthsfwd = 0.1 xjbvs = 1 bvs = 12.69
+ jss = 2.1483E-5 jsws = 4.02E-12 cjs = {sw_psd_nw_cj}
+ mjs = 0.33956 mjsws = 0.24676 cjsws = {9.960545E-11*sw_func_psd_nw_cj}
+ cjswgs = {1.47314E-10*sw_func_psd_nw_cj} mjswgs = 0.81 pbs = 0.6587
+ pbsws = 1 pbswgs = 3 xrcrg1 = 12
+ xrcrg2 = 1 rbpb = 50 rbpd = 50
+ rbps = 50 rbdb = 50 rbsb = 50
+ gbmin = 1E-12 tnom = 30 ute = -2.39937
+ lute = 4.509132E-7 wute = 5.515497E-7 pute = -1.950764E-13
+ kt1 = -0.882734 lkt1 = 1.228087E-7 wkt1 = 2.402451E-8
+ pkt1 = -1.814664E-14 kt1l = 0 kt2 = -0.019032
+ ua1 = 5.52E-10 ub1 = -7.043152E-18 lub1 = 1.551534E-24
+ wub1 = 6.205801E-24 pub1 = -2.103801E-30 uc1 = -8.475202E-12
+ wuc1 = -9.82516E-17 at = 3.937727E3 lat = 9.148196E-3
+ wat = 4.18415E-2 pat = -2.721996E-8 prt = 0
+ njs = 1.3632 xtis = 10 tpb = 1.671E-3
+ tpbsw = 0 tpbswg = 0 tcj = 9.6E-4
+ tcjsw = 3E-5 tcjswg = 0 tvoff = 0
+ tvfbsdoff = 0 saref = 2.02E-6 sbref = 2.01E-6
+ wlod = 0 ku0 = 7E-8 kvsat = 0.4
+ kvth0 = 3.5E-8 tku0 = 0 llodku0 = 0
+ wlodku0 = 1 llodvth = 0 wlodvth = 1
+ lku0 = 0 wku0 = 0 pku0 = 0
+ lkvth0 = 0 wkvth0 = 6.5E-7 pkvth0 = 0
+ stk2 = 0 lodk2 = 1 steta0 = 0
+ lodeta0 = 1

.model phv_model.36 pmos
+ level = 54 lmin = 8E-6 lmax = 2.02E-5 wmin = 7.5E-7
+ wmax = 1E-6 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 1.175E-8
+ toxm = 1.175E-8 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 1E23 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {1.2277E-8+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {4.5375E-8-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = -4.7338E-9 dwb = 0 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = -0.960189 k1 = 0.58485
+ k2 = 2.52294E-2 k3 = -2.2405 k3b = -0.172
+ w0 = 0 lpe0 = 0 lpeb = 0
+ vbm = -3 dvtp0 = 0 dvtp1 = 0
+ dvt0 = 4.657 dvt1 = 0.34864 dvt2 = -0.030206
+ dvt0w = -2.2 dvt1w = 1.0163E6 dvt2w = 0
+ vfbsdoff = 0 u0 = 1.86026E-2 ua = 2.250479E-9
+ ub = 2.47633E-19 uc = -4.510858E-11 ud = 0
+ up = 0 lp = 1 eu = 1.67
+ vsat = 8.0156E4 a0 = 0.906425 ags = 0.137596
+ b0 = 0 b1 = 0 keta = -8.1819E-3
+ a1 = 0 a2 = 0.5 rdsw = 788.47
+ rdswmin = 0 rdw = 0 rdwmin = 0
+ rsw = 0 rswmin = 0 prwb = 0.053538
+ prwg = 0 wr = 1 voff = -0.10768
+ voffl = 0 minv = 0 nfactor = 1.59862
+ eta0 = 0.08 etab = -0.07 dsub = 0.56
+ cit = 5E-6 cdsc = 0 cdscb = 0
+ cdscd = 0 pclm = 8.35312E-2 pdiblc1 = 0.39
+ pdiblc2 = 3.438067E-3 pdiblcb = -0.025 drout = 0.56
+ pscbe1 = 2.247176E8 pscbe2 = 1.499872E-8 pvag = 0
+ delta = 0.01 fprout = 0 pdits = 0
+ pditsl = 0 pditsd = 0 lambda = 0
+ vtl = 0 lc = 5E-9 xn = 3
+ alpha0 = 6.424264E-5 alpha1 = 0 beta0 = 39.039478
+ aigbacc = 0.43 bigbacc = 0.054 cigbacc = 0.075
+ nigbacc = 1 aigbinv = 0.35 bigbinv = 0.03
+ cigbinv = 6E-3 eigbinv = 1.1 nigbinv = 3
+ aigc = 0.43 bigc = 0.054 cigc = 0.075
+ aigsd = 0.43 bigsd = 0.054 cigsd = 0.075
+ dlcig = 0 nigc = 1 poxedge = 1
+ pigcd = 1 ntox = 1 toxref = 1.175E-8
+ agidl = 2E-8 bgidl = 1.5204E9 cgidl = 1.4E3
+ egidl = 1.519935 noia = 3E40 noib = 8.53E24
+ noic = 8.4E7 em = 4.1E7 af = 1
+ ef = 0.88 kf = 0 lintnoi = 0
+ tnoia = 1.5 tnoib = 3.5 ntnoi = 1
+ rnoia = 0.577 rnoib = 0.37 xpart = 0
+ cgso = {1.94171E-10/sw_func_tox_hv_ratio} cgdo = {1.94171E-10/sw_func_tox_hv_ratio} cgbo = {0/sw_func_tox_hv_ratio}
+ ckappas = 0.6 cf = 1.2E-11 clc = 1E-7
+ cle = 0.6 dlc = 4.4983E-8 dwc = 0
+ vfbcv = -0.144689 noff = 4 voffcv = 0
+ acde = 0.401 moin = 15.773 cgsl = {9.82591E-12/sw_func_tox_hv_ratio}
+ cgdl = {9.82591E-12/sw_func_tox_hv_ratio} ijthsrev = 0.1 ijthsfwd = 0.1
+ xjbvs = 1 bvs = 12.69 jss = 2.1483E-5
+ jsws = 4.02E-12 cjs = {sw_psd_nw_cj} mjs = 0.33956
+ mjsws = 0.24676 cjsws = {9.960545E-11*sw_func_psd_nw_cj} cjswgs = {1.47314E-10*sw_func_psd_nw_cj}
+ mjswgs = 0.81 pbs = 0.6587 pbsws = 1
+ pbswgs = 3 xrcrg1 = 12 xrcrg2 = 1
+ rbpb = 50 rbpd = 50 rbps = 50
+ rbdb = 50 rbsb = 50 gbmin = 1E-12
+ tnom = 30 ute = -1.5561 kt1 = -0.556
+ kt1l = 0 kt2 = -0.019032 ua1 = 2.2096E-11
+ ub1 = -3.0767E-18 uc1 = -1.092E-10 at = 1.5109E5
+ prt = 0 njs = 1.3632 xtis = 10
+ tpb = 1.671E-3 tpbsw = 0 tpbswg = 0
+ tcj = 9.6E-4 tcjsw = 3E-5 tcjswg = 0
+ tvoff = 0 tvfbsdoff = 0 saref = 3E-6
+ sbref = 3E-6 wlod = 0 ku0 = 7E-8
+ kvsat = 0.4 kvth0 = 3.5E-8 tku0 = 0
+ llodku0 = 0 wlodku0 = 1 llodvth = 0
+ wlodvth = 1 lku0 = 0 wku0 = 0
+ pku0 = 0 lkvth0 = 0 wkvth0 = 6.5E-7
+ pkvth0 = 0 stk2 = 0 lodk2 = 1
+ steta0 = 0 lodeta0 = 1

.model phv_model.37 pmos
+ level = 54 lmin = 4E-6 lmax = 8E-6 wmin = 7.5E-7
+ wmax = 1E-6 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 1.175E-8
+ toxm = 1.175E-8 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 1E23 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {1.2277E-8+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {4.5375E-8-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = -4.7338E-9 dwb = 0 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = -0.973912 lvth0 = 1.08542E-7
+ k1 = 0.565059 lk1 = 1.565286E-7 k2 = 3.14423E-2
+ lk2 = -4.913982E-8 k3 = -2.2405 k3b = -0.172
+ w0 = 0 lpe0 = 0 lpeb = 0
+ vbm = -3 dvtp0 = 0 dvtp1 = 0
+ dvt0 = 4.657 dvt1 = 0.34864 dvt2 = -0.030206
+ dvt0w = -2.2 dvt1w = 1.0163E6 dvt2w = 0
+ vfbsdoff = 0 u0 = 1.93395E-2 lu0 = -5.82843E-9
+ ua = 2.527816E-9 lua = -2.193531E-15 ub = 1.196569E-19
+ lub = 1.012195E-24 uc = -5.99701E-11 luc = 1.175435E-16
+ ud = 0 up = 0 lp = 1
+ eu = 1.67 vsat = 4.099118E4 lvsat = 0.309764
+ a0 = 0.944463 la0 = -3.008469E-7 ags = 0.137255
+ lags = 2.698554E-9 b0 = 0 b1 = 0
+ keta = -6.573928E-3 lketa = -1.271785E-8 a1 = 0
+ a2 = 0.5 rdsw = 788.47 rdswmin = 0
+ rdw = 0 rdwmin = 0 rsw = 0
+ rswmin = 0 prwb = 0.053538 prwg = 0
+ wr = 1 voff = -0.118049 lvoff = 8.201056E-8
+ voffl = 0 minv = 0 nfactor = 1.538633
+ lnfactor = 4.744557E-7 eta0 = 0.08 etab = -0.07
+ dsub = 0.56 cit = 1.134375E-7 lcit = 3.864904E-11
+ cdsc = 0 cdscb = 0 cdscd = 0
+ pclm = -0.727727 lpclm = 6.416446E-6 pdiblc1 = 0.39
+ pdiblc2 = 5.537399E-3 lpdiblc2 = -1.660414E-8 pdiblcb = -0.025
+ drout = 0.56 pscbe1 = 2.243843E8 lpscbe1 = 2.636329
+ pscbe2 = 1.499872E-8 pvag = 0 delta = 0.01
+ fprout = 0 pdits = 0 pditsl = 0
+ pditsd = 0 lambda = 0 vtl = 0
+ lc = 5E-9 xn = 3 alpha0 = 1.270277E-4
+ lalpha0 = -4.965826E-10 alpha1 = -9.773125E-11 lalpha1 = 7.729809E-16
+ beta0 = 74.26131 lbeta0 = -2.785783E-4 aigbacc = 0.43
+ bigbacc = 0.054 cigbacc = 0.075 nigbacc = 1
+ aigbinv = 0.35 bigbinv = 0.03 cigbinv = 6E-3
+ eigbinv = 1.1 nigbinv = 3 aigc = 0.43
+ bigc = 0.054 cigc = 0.075 aigsd = 0.43
+ bigsd = 0.054 cigsd = 0.075 dlcig = 0
+ nigc = 1 poxedge = 1 pigcd = 1
+ ntox = 1 toxref = 1.175E-8 agidl = 6.70855E-9
+ lagidl = 1.051254E-13 bgidl = 1.567409E9 lbgidl = -371.803808
+ cgidl = 2.2874E3 lcgidl = -7.018666E-3 egidl = 1.050762
+ legidl = 3.710809E-6 noia = 3E40 noib = 8.53E24
+ noic = 8.4E7 em = 4.1E7 af = 1
+ ef = 0.88 kf = 0 lintnoi = 0
+ tnoia = 1.5 tnoib = 3.5 ntnoi = 1
+ rnoia = 0.577 rnoib = 0.37 xpart = 0
+ cgso = {1.94171E-10/sw_func_tox_hv_ratio} cgdo = {1.94171E-10/sw_func_tox_hv_ratio} cgbo = {0/sw_func_tox_hv_ratio}
+ ckappas = 0.6 cf = 1.2E-11 clc = 1E-7
+ cle = 0.6 dlc = 4.4983E-8 dwc = 0
+ vfbcv = -0.144689 noff = 4 voffcv = 0
+ acde = 0.401 moin = 15.773 cgsl = {9.82591E-12/sw_func_tox_hv_ratio}
+ cgdl = {9.82591E-12/sw_func_tox_hv_ratio} ijthsrev = 0.1 ijthsfwd = 0.1
+ xjbvs = 1 bvs = 12.69 jss = 2.1483E-5
+ jsws = 4.02E-12 cjs = {sw_psd_nw_cj} mjs = 0.33956
+ mjsws = 0.24676 cjsws = {9.960545E-11*sw_func_psd_nw_cj} cjswgs = {1.47314E-10*sw_func_psd_nw_cj}
+ mjswgs = 0.81 pbs = 0.6587 pbsws = 1
+ pbswgs = 3 xrcrg1 = 12 xrcrg2 = 1
+ rbpb = 50 rbpd = 50 rbps = 50
+ rbdb = 50 rbsb = 50 gbmin = 1E-12
+ tnom = 30 ute = -1.698494 lute = 1.126233E-6
+ kt1 = -0.536454 lkt1 = -1.545962E-7 kt1l = 0
+ kt2 = -0.019032 ua1 = 2.2096E-11 ub1 = -3.738243E-18
+ lub1 = 5.232308E-24 uc1 = -1.092E-10 at = 8.408545E4
+ lat = 0.529956 prt = 0 njs = 1.3632
+ xtis = 10 tpb = 1.671E-3 tpbsw = 0
+ tpbswg = 0 tcj = 9.6E-4 tcjsw = 3E-5
+ tcjswg = 0 tvoff = 0 tvfbsdoff = 0
+ saref = 3E-6 sbref = 3E-6 wlod = 0
+ ku0 = 7E-8 kvsat = 0.4 kvth0 = 3.5E-8
+ tku0 = 0 llodku0 = 0 wlodku0 = 1
+ llodvth = 0 wlodvth = 1 lku0 = 0
+ wku0 = 0 pku0 = 0 lkvth0 = 0
+ wkvth0 = 6.5E-7 pkvth0 = 0 stk2 = 0
+ lodk2 = 1 steta0 = 0 lodeta0 = 1

.model phv_model.38 pmos
+ level = 54 lmin = 2E-6 lmax = 4E-6 wmin = 7.5E-7
+ wmax = 1E-6 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 1.175E-8
+ toxm = 1.175E-8 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 1E23 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {1.2277E-8+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {4.5375E-8-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = -4.7338E-9 dwb = 0 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = -0.911019 lvth0 = -1.373232E-7
+ wvth0 = -4.356106E-8 pvth0 = 1.702911E-13 k1 = 0.523006
+ lk1 = 3.209258E-7 wk1 = 9.089858E-8 pk1 = -3.553453E-13
+ k2 = 4.09019E-2 lk2 = -8.611959E-8 wk2 = -2.699186E-8
+ pk2 = 1.055179E-13 k3 = -2.2405 k3b = -0.172
+ w0 = 0 lpe0 = 0 lpeb = 0
+ vbm = -3 dvtp0 = 0 dvtp1 = 0
+ dvt0 = 4.657 dvt1 = 0.34864 dvt2 = -0.030206
+ dvt0w = -2.2 dvt1w = 1.0163E6 dvt2w = 0
+ vfbsdoff = 0 u0 = 1.88578E-2 lu0 = -3.94534E-9
+ wu0 = -1.399687E-10 pu0 = 5.471726E-16 ua = 3.319929E-9
+ lua = -5.290096E-15 wua = -1.026412E-15 pua = 4.012501E-21
+ ub = -2.126939E-18 lub = 9.794701E-24 wub = 2.256765E-24
+ pub = -8.82226E-30 uc = -2.031571E-11 luc = -3.747544E-17
+ wuc = -2.572542E-17 puc = 1.005671E-22 ud = 0
+ up = 0 lp = 1 eu = 1.67
+ vsat = 2.623576E5 lvsat = -0.555612 wvsat = -4.62977E-2
+ pvsat = 1.809895E-7 a0 = 0.217973 la0 = 2.539184E-6
+ wa0 = 5.599585E-7 pa0 = -2.189018E-12 ags = -1.132622
+ lags = 4.966965E-6 wags = 7.177946E-7 pags = -2.806038E-12
+ b0 = 1.847916E-7 lb0 = -7.223967E-13 wb0 = -1.802543E-13
+ pb0 = 7.04659E-19 b1 = 1.080622E-9 lb1 = -4.224422E-15
+ wb1 = -1.054088E-15 pb1 = 4.120695E-21 keta = 0.305672
+ lketa = -1.233365E-6 wketa = -2.099287E-7 pketa = 8.206638E-13
+ a1 = 0 a2 = 0.5 rdsw = 788.47
+ rdswmin = 0 rdw = 0 rdwmin = 0
+ rsw = 0 rswmin = 0 prwb = 0.053538
+ prwg = 0 wr = 1 voff = -7.86139E-2
+ lvoff = -7.215155E-8 wvoff = -2.816533E-8 pvoff = 1.101053E-13
+ voffl = 0 minv = 0 nfactor = 2.122423
+ lnfactor = -1.807729E-6 wnfactor = -4.714621E-7 pnfactor = 1.843063E-12
+ eta0 = 0.322577 leta0 = -9.482939E-7 weta0 = -1.621259E-7
+ peta0 = 6.337906E-13 etab = -0.13441 letab = 2.517953E-7
+ wetab = -1.75096E-9 petab = 6.844939E-15 dsub = 1.001391
+ ldsub = -1.725509E-6 wdsub = -1.511978E-7 pdsub = 5.910701E-13
+ cit = 2.137543E-5 lcit = -4.446941E-11 wcit = -8.252263E-12
+ pcit = 3.226016E-17 cdsc = 0 cdscb = 0
+ cdscd = 0 pclm = -2.061244 lpclm = 1.16295E-5
+ wpclm = 1.98003E-6 ppclm = -7.740432E-12 pdiblc1 = 0.820472
+ lpdiblc1 = -1.682822E-6 wpdiblc1 = -4.207478E-7 ppdiblc1 = 1.644808E-12
+ pdiblc2 = 3.341699E-3 lpdiblc2 = -8.020604E-9 wpdiblc2 = -2.001321E-9
+ ppdiblc2 = 7.823666E-15 pdiblcb = -0.025 drout = -0.102165
+ ldrout = 2.588568E-6 wdrout = 5.732735E-7 pdrout = -2.241069E-12
+ pscbe1 = 5.606935E7 lpscbe1 = 660.621495 wpscbe1 = 85.83466
+ ppscbe1 = -3.355491E-4 pscbe2 = 1.453255E-8 lpscbe2 = 1.856278E-15
+ wpscbe2 = 6.861816E-16 ppscbe2 = -2.682455E-21 pvag = 0
+ delta = 0.01 fprout = 0 pdits = 0
+ pditsl = 0 pditsd = 0 lambda = 0
+ vtl = 0 lc = 5E-9 xn = 3
+ alpha0 = -1.19105E-3 lalpha0 = 4.656113E-9 walpha0 = 8.640426E-10
+ palpha0 = -3.377759E-15 alpha1 = 4.724741E-10 lalpha1 = -1.456094E-15
+ walpha1 = -2.702098E-16 palpha1 = 1.056318E-21 beta0 = -191.966106
+ lbeta0 = 7.621712E-4 wbeta0 = 1.414374E-4 pbeta0 = -5.529141E-10
+ aigbacc = 0.43 bigbacc = 0.054 cigbacc = 0.075
+ nigbacc = 1 aigbinv = 0.35 bigbinv = 0.03
+ cigbinv = 6E-3 eigbinv = 1.1 nigbinv = 3
+ aigc = 0.43 bigc = 0.054 cigc = 0.075
+ aigsd = 0.43 bigsd = 0.054 cigsd = 0.075
+ dlcig = 0 nigc = 1 poxedge = 1
+ pigcd = 1 ntox = 1 toxref = 1.175E-8
+ agidl = -8.30217E-8 lagidl = 4.559034E-13 wagidl = 1.077986E-13
+ pagidl = -4.214116E-19 bgidl = -2.535852E8 lbgidl = 6.746917E3
+ wbgidl = 1.559381E3 pbgidl = -6.09601E-3 cgidl = 2.458986E3
+ lcgidl = -7.689442E-3 wcgidl = -2.242741E-3 pcgidl = 8.767437E-9
+ egidl = 1.001943 legidl = 3.901654E-6 wegidl = 1.479119E-6
+ pegidl = -5.782244E-12 noia = 3E40 noib = 8.53E24
+ noic = 8.4E7 em = 4.1E7 af = 1
+ ef = 0.88 kf = 0 lintnoi = 0
+ tnoia = 1.5 tnoib = 3.5 ntnoi = 1
+ rnoia = 0.577 rnoib = 0.37 xpart = 0
+ cgso = {1.94171E-10/sw_func_tox_hv_ratio} cgdo = {1.94171E-10/sw_func_tox_hv_ratio} cgbo = {0/sw_func_tox_hv_ratio}
+ ckappas = 0.6 cf = 1.2E-11 clc = 1E-7
+ cle = 0.6 dlc = 4.4983E-8 dwc = 0
+ vfbcv = -0.144689 noff = 4 voffcv = 0
+ acde = 0.401 moin = 15.773 cgsl = {9.82591E-12/sw_func_tox_hv_ratio}
+ cgdl = {9.82591E-12/sw_func_tox_hv_ratio} ijthsrev = 0.1 ijthsfwd = 0.1
+ xjbvs = 1 bvs = 12.69 jss = 2.1483E-5
+ jsws = 4.02E-12 cjs = {sw_psd_nw_cj} mjs = 0.33956
+ mjsws = 0.24676 cjsws = {9.960545E-11*sw_func_psd_nw_cj} cjswgs = {1.47314E-10*sw_func_psd_nw_cj}
+ mjswgs = 0.81 pbs = 0.6587 pbsws = 1
+ pbswgs = 3 xrcrg1 = 12 xrcrg2 = 1
+ rbpb = 50 rbpd = 50 rbps = 50
+ rbdb = 50 rbsb = 50 gbmin = 1E-12
+ tnom = 30 ute = -1.544126 lute = 5.227677E-7
+ wute = 1.242965E-7 pute = -4.859061E-13 kt1 = -0.630183
+ lkt1 = 2.118166E-7 wkt1 = 8.916924E-8 pkt1 = -3.485848E-13
+ kt1l = 0 kt2 = -0.019032 ua1 = -1.307164E-9
+ lua1 = 5.19641E-15 wua1 = 5.970556E-16 pua1 = -2.33404E-21
+ ub1 = -4.205291E-18 lub1 = 7.058116E-24 wub1 = 2.134658E-24
+ pub1 = -8.34491E-30 uc1 = -1.092E-10 at = 4.630237E5
+ lat = -0.951409 wat = -4.85405E-2 pat = 1.897569E-7
+ prt = 0 njs = 1.3632 xtis = 10
+ tpb = 1.671E-3 tpbsw = 0 tpbswg = 0
+ tcj = 9.6E-4 tcjsw = 3E-5 tcjswg = 0
+ tvoff = 0 tvfbsdoff = 0 saref = 3E-6
+ sbref = 3E-6 wlod = 0 ku0 = 7E-8
+ kvsat = 0.4 kvth0 = 3.5E-8 tku0 = 0
+ llodku0 = 0 wlodku0 = 1 llodvth = 0
+ wlodvth = 1 lku0 = 0 wku0 = 0
+ pku0 = 0 lkvth0 = 0 wkvth0 = 6.5E-7
+ pkvth0 = 0 stk2 = 0 lodk2 = 1
+ steta0 = 0 lodeta0 = 1

.model phv_model.39 pmos
+ level = 54 lmin = 1E-6 lmax = 2E-6 wmin = 7.5E-7
+ wmax = 1E-6 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 1.175E-8
+ toxm = 1.175E-8 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 1E23 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {1.2277E-8+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {4.5375E-8-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = -4.7338E-9 dwb = 0 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = -1.017332 lvth0 = 6.56536E-8
+ wvth0 = 6.283705E-8 pvth0 = -3.28495E-14 k1 = 0.681198
+ lk1 = 1.88979E-8 wk1 = -8.803863E-8 pk1 = -1.370941E-14
+ k2 = -3.424217E-3 lk2 = -1.49002E-9 wk2 = 2.742596E-8
+ pk2 = 1.620693E-15 k3 = -2.2405 k3b = -0.172
+ w0 = 0 lpe0 = 0 lpeb = 0
+ vbm = -3 dvtp0 = 0 dvtp1 = 0
+ dvt0 = 4.657 dvt1 = 0.34864 dvt2 = -0.030206
+ dvt0w = -2.2 dvt1w = 1.0163E6 dvt2w = 0
+ vfbsdoff = 0 u0 = 2.31231E-2 lu0 = -1.208875E-8
+ wu0 = -4.315801E-9 pu0 = 8.51988E-15 ua = 3.089014E-9
+ lua = -4.849222E-15 wua = -7.672382E-16 pua = 3.517673E-21
+ ub = 7.794534E-19 lub = 4.245671E-24 wub = -7.737929E-25
+ pub = -3.036167E-30 uc = -7.576028E-11 luc = 6.838209E-17
+ wuc = 5.293091E-17 puc = -4.960752E-23 ud = 0
+ up = 0 lp = 1 eu = 1.67
+ vsat = -3.41136E4 lvsat = 1.04253E-2 wvsat = 3.17953E-2
+ pvsat = 3.189034E-8 a0 = 1.807298 la0 = -4.95235E-7
+ wa0 = -7.747457E-7 pa0 = 3.592662E-13 ags = 1.446656
+ lags = 4.247965E-8 wags = -7.357719E-7 pags = -3.081669E-14
+ b0 = -1.322576E-7 lb0 = -1.170705E-13 wb0 = 1.290101E-13
+ pb0 = 1.141959E-19 b1 = 5.695486E-10 lb1 = -3.248655E-15
+ wb1 = -5.555639E-16 pb1 = 3.168887E-21 keta = -0.425643
+ lketa = 1.628978E-7 wketa = 2.787898E-7 pketa = -1.12422E-13
+ a1 = 0 a2 = 0.5 rdsw = 788.47
+ rdswmin = 0 rdw = 0 rdwmin = 0
+ rsw = 0 rswmin = 0 prwb = 0.053538
+ prwg = 0 wr = 1 voff = -0.13951
+ lvoff = 4.41152E-8 wvoff = 4.626626E-8 pvoff = -3.200319E-14
+ voffl = 0 minv = 0 nfactor = 1.040807
+ lnfactor = 2.573468E-7 wnfactor = 6.719947E-7 pnfactor = -3.400817E-13
+ eta0 = -0.37742 leta0 = 3.881752E-7 weta0 = 3.33082E-7
+ peta0 = -3.116851E-13 etab = -1.34909E-2 letab = 2.093026E-8
+ wetab = 1.265011E-8 petab = -2.06503E-14 dsub = -7.23543E-2
+ ldsub = 3.245399E-7 wdsub = 2.816979E-7 pdsub = -2.354361E-13
+ cit = 4.987618E-6 lcit = -1.318098E-11 wcit = 3.636212E-12
+ pcit = 9.562087E-18 cdsc = 0 cdscb = 0
+ cdscd = 0 pclm = 6.284773 lpclm = -4.305137E-6
+ wpclm = -3.709941E-6 ppclm = 3.123144E-12 pdiblc1 = 0.172007
+ lpdiblc1 = -4.447397E-7 wpdiblc1 = 2.717617E-7 ppdiblc1 = 3.226346E-13
+ pdiblc2 = -3.423145E-3 lpdiblc2 = 4.895175E-9 wpdiblc2 = 3.956437E-9
+ ppdiblc2 = -3.551185E-15 pdiblcb = -0.025 drout = -3.06259E-2
+ ldrout = 2.451982E-6 wdrout = 3.311424E-7 pdrout = -1.778781E-12
+ pscbe1 = 3.980557E8 lpscbe1 = 7.683994 wpscbe1 = -86.994892
+ ppscbe1 = -5.574323E-6 pscbe2 = 1.674477E-8 lpscbe2 = -2.367412E-15
+ wpscbe2 = -1.618328E-15 ppscbe2 = 1.71743E-21 pvag = 0
+ delta = 0.01 fprout = 0 pdits = 0
+ pditsl = 0 pditsd = 0 lambda = 0
+ vtl = 0 lc = 5E-9 xn = 3
+ alpha0 = 2.118745E-3 lalpha0 = -1.663114E-9 walpha0 = -1.537035E-9
+ palpha0 = 1.206499E-15 alpha1 = -2.901784E-10 walpha1 = 2.830534E-16
+ beta0 = 226.361681 lbeta0 = -3.652108E-5 wbeta0 = -1.620368E-4
+ pbeta0 = 2.649407E-11 aigbacc = 0.43 bigbacc = 0.054
+ cigbacc = 0.075 nigbacc = 1 aigbinv = 0.35
+ bigbinv = 0.03 cigbinv = 6E-3 eigbinv = 1.1
+ nigbinv = 3 aigc = 0.43 bigc = 0.054
+ cigc = 0.075 aigsd = 0.43 bigsd = 0.054
+ cigsd = 0.075 dlcig = 0 nigc = 1
+ poxedge = 1 pigcd = 1 ntox = 1
+ toxref = 1.175E-8 agidl = 2.909975E-7 lagidl = -2.581927E-13
+ wagidl = -2.110263E-13 pagidl = 1.873049E-19 bgidl = 3.502305E9
+ lbgidl = -424.017387 wbgidl = -1.794612E3 pbgidl = 3.076017E-4
+ cgidl = -1.649657E3 lcgidl = 1.549851E-4 wcgidl = 2.85409E-3
+ pcgidl = -9.636877E-10 egidl = 7.859971 legidl = -9.192036E-6
+ wegidl = -5.042065E-6 pegidl = 6.668326E-12 noia = 3E40
+ noib = 8.53E24 noic = 8.4E7 em = 4.1E7
+ af = 1 ef = 0.88 kf = 0
+ lintnoi = 0 tnoia = 1.5 tnoib = 3.5
+ ntnoi = 1 rnoia = 0.577 rnoib = 0.37
+ xpart = 0 cgso = {1.94171E-10/sw_func_tox_hv_ratio} cgdo = {1.94171E-10/sw_func_tox_hv_ratio}
+ cgbo = {0/sw_func_tox_hv_ratio} ckappas = 0.6 cf = 1.2E-11
+ clc = 1E-7 cle = 0.6 dlc = 4.4983E-8
+ dwc = 0 vfbcv = -0.144689 noff = 4
+ voffcv = 0 acde = 0.401 moin = 15.773
+ cgsl = {9.82591E-12/sw_func_tox_hv_ratio} cgdl = {9.82591E-12/sw_func_tox_hv_ratio} ijthsrev = 0.1
+ ijthsfwd = 0.1 xjbvs = 1 bvs = 12.69
+ jss = 2.1483E-5 jsws = 4.02E-12 cjs = {sw_psd_nw_cj}
+ mjs = 0.33956 mjsws = 0.24676 cjsws = {9.960545E-11*sw_func_psd_nw_cj}
+ cjswgs = {1.47314E-10*sw_func_psd_nw_cj} mjswgs = 0.81 pbs = 0.6587
+ pbsws = 1 pbswgs = 3 xrcrg1 = 12
+ xrcrg2 = 1 rbpb = 50 rbpd = 50
+ rbps = 50 rbdb = 50 rbsb = 50
+ gbmin = 1E-12 tnom = 30 ute = -1.107124
+ lute = -3.115783E-7 wute = -2.48593E-7 pute = 2.260332E-13
+ kt1 = -0.437644 lkt1 = -1.557891E-7 wkt1 = -1.526019E-7
+ pkt1 = 1.130166E-13 kt1l = 0 kt2 = -0.019032
+ ua1 = 2.198437E-9 lua1 = -1.496659E-15 wua1 = -1.194111E-15
+ pua1 = 1.085746E-21 ub1 = 2.29419E-18 lub1 = -5.351018E-24
+ wub1 = -4.269315E-24 pub1 = 3.881875E-30 uc1 = -1.092E-10
+ at = -9.465808E4 lat = 0.113345 wat = 0.097081
+ pat = -8.827088E-8 prt = 0 njs = 1.3632
+ xtis = 10 tpb = 1.671E-3 tpbsw = 0
+ tpbswg = 0 tcj = 9.6E-4 tcjsw = 3E-5
+ tcjswg = 0 tvoff = 0 tvfbsdoff = 0
+ saref = 3E-6 sbref = 3E-6 wlod = 0
+ ku0 = 7E-8 kvsat = 0.4 kvth0 = 3.5E-8
+ tku0 = 0 llodku0 = 0 wlodku0 = 1
+ llodvth = 0 wlodvth = 1 lku0 = 0
+ wku0 = 0 pku0 = 0 lkvth0 = 0
+ wkvth0 = 6.5E-7 pkvth0 = 0 stk2 = 0
+ lodk2 = 1 steta0 = 0 lodeta0 = 1

.model phv_model.40 pmos
+ level = 54 lmin = 8E-7 lmax = 1E-6 wmin = 7.5E-7
+ wmax = 1E-6 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 1.175E-8
+ toxm = 1.175E-8 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 1E23 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {1.2277E-8+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {4.5375E-8-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = -4.7338E-9 dwb = 0 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = -0.880397 lvth0 = -5.885439E-8
+ wvth0 = -2.483508E-8 pvth0 = 4.686638E-14 k1 = 0.969169
+ lk1 = -2.429395E-7 wk1 = -2.969459E-7 pk1 = 1.762395E-13
+ k2 = -8.62169E-2 lk2 = 7.378921E-8 wk2 = 8.099777E-8
+ pk2 = -4.708948E-14 k3 = -2.2405 k3b = -0.172
+ w0 = 0 lpe0 = 0 lpeb = 0
+ vbm = -3 dvtp0 = 0 dvtp1 = 0
+ dvt0 = 4.657 dvt1 = 0.34864 dvt2 = -0.030206
+ dvt0w = -2.2 dvt1w = 1.0163E6 dvt2w = 0
+ vfbsdoff = 0 u0 = -4.306541E-3 lu0 = 1.285161E-8
+ wu0 = 1.586893E-8 pu0 = -9.833087E-15 ua = -8.401167E-9
+ lua = 5.598225E-15 wua = 7.563272E-15 pua = -4.056843E-21
+ ub = 1.080191E-17 lub = -4.867248E-24 wub = -7.939193E-24
+ pub = 3.478973E-30 uc = -5.147071E-12 luc = 4.177037E-18
+ wuc = 1.704847E-18 puc = -3.030215E-24 ud = 0
+ up = 0 lp = 1 eu = 1.67
+ vsat = -1.43688E5 lvsat = 0.110056 wvsat = 0.147108
+ pvsat = -7.295731E-8 a0 = 2.334242 la0 = -9.743593E-7
+ wa0 = -1.157016E-6 pa0 = 7.068451E-13 ags = 1.058912
+ lags = 3.950353E-7 wags = -4.54485E-7 pags = -2.865768E-13
+ b0 = -1.186628E-6 lb0 = 8.416162E-13 wb0 = 1.157492E-12
+ pb0 = -8.209511E-19 b1 = -1.365396E-8 lb1 = 9.684074E-15
+ wb1 = 1.33187E-14 pb1 = -9.446291E-21 keta = -0.562199
+ lketa = 2.870612E-7 wketa = 3.841792E-7 pketa = -2.082474E-13
+ a1 = 0 a2 = 0.5 rdsw = 788.47
+ rdswmin = 0 rdw = 0 rdwmin = 0
+ rsw = 0 rswmin = 0 prwb = 0.053538
+ prwg = 0 wr = 1 voff = -3.60546E-2
+ lvoff = -4.995202E-8 wvoff = -2.878537E-8 pvoff = 3.62375E-14
+ voffl = 0 minv = 0 nfactor = 2.002304
+ lnfactor = -6.168942E-7 wnfactor = -1.85138E-7 pnfactor = 4.392662E-13
+ eta0 = 0.502204 leta0 = -4.116233E-7 weta0 = -3.381256E-7
+ peta0 = 2.986105E-13 etab = 5.53049E-2 letab = -4.162229E-8
+ wetab = -4.326963E-8 petab = 3.019473E-14 dsub = 0.875512
+ ldsub = -5.373073E-7 wdsub = -4.059277E-7 pdsub = 3.897875E-13
+ cit = -7.869243E-5 lcit = 6.29051E-11 wcit = 6.434157E-11
+ pcit = -4.563426E-17 cdsc = 0 cdscb = 0
+ cdscd = 0 pclm = 3.144811 lpclm = -1.450126E-6
+ wpclm = -1.432068E-6 ppclm = 1.051988E-12 pdiblc1 = -2.100465
+ lpdiblc1 = 1.621505E-6 wpdiblc1 = 1.920317E-6 ppdiblc1 = -1.176314E-12
+ pdiblc2 = -0.061562 lpdiblc2 = 5.775794E-8 wpdiblc2 = 4.613305E-8
+ ppdiblc2 = -4.190027E-14 pdiblcb = -0.025 drout = 8.946579
+ ldrout = -5.710542E-6 wdrout = -6.181335E-6 pdrout = 4.14269E-12
+ pscbe1 = -3.944036E8 lpscbe1 = 728.227607 wpscbe1 = 487.891533
+ ppscbe1 = -5.282898E-4 pscbe2 = 2.706508E-8 lpscbe2 = -1.175115E-14
+ wpscbe2 = -9.105154E-15 ppscbe2 = 8.524826E-21 pvag = 0
+ delta = 0.01 fprout = 0 pdits = 0
+ pditsl = 0 pditsd = 0 lambda = 0
+ vtl = 0 lc = 5E-9 xn = 3
+ alpha0 = 8.676986E-4 lalpha0 = -5.255995E-10 walpha0 = -6.294684E-10
+ palpha0 = 3.812941E-16 alpha1 = -2.901784E-10 walpha1 = 2.830534E-16
+ beta0 = 220.844424 lbeta0 = -3.150451E-5 wbeta0 = -1.580344E-4
+ pbeta0 = 2.285482E-11 aigbacc = 0.43 bigbacc = 0.054
+ cigbacc = 0.075 nigbacc = 1 aigbinv = 0.35
+ bigbinv = 0.03 cigbinv = 6E-3 eigbinv = 1.1
+ nigbinv = 3 aigc = 0.43 bigc = 0.054
+ cigc = 0.075 aigsd = 0.43 bigsd = 0.054
+ cigsd = 0.075 dlcig = 0 nigc = 1
+ poxedge = 1 pigcd = 1 ntox = 1
+ toxref = 1.175E-8 agidl = -7.285304E-8 lagidl = 7.263836E-14
+ wagidl = 5.25818E-14 pagidl = -5.238082E-20 bgidl = -3.62326E8
+ lbgidl = 3.089899E3 wbgidl = 1.008969E3 pbgidl = -2.241555E-3
+ cgidl = -3.552217E3 lcgidl = 1.884889E-3 wcgidl = 3.298079E-3
+ pcgidl = -1.367385E-9 egidl = -3.10899 legidl = 7.814916E-7
+ wegidl = 2.915323E-6 pegidl = -5.6693E-13 noia = 3E40
+ noib = 8.53E24 noic = 8.4E7 em = 4.1E7
+ af = 1 ef = 0.88 kf = 0
+ lintnoi = 0 tnoia = 1.5 tnoib = 3.5
+ ntnoi = 1 rnoia = 0.577 rnoib = 0.37
+ xpart = 0 cgso = {1.94171E-10/sw_func_tox_hv_ratio} cgdo = {1.94171E-10/sw_func_tox_hv_ratio}
+ cgbo = {0/sw_func_tox_hv_ratio} ckappas = 0.6 cf = 1.2E-11
+ clc = 1E-7 cle = 0.6 dlc = 4.4983E-8
+ dwc = 0 vfbcv = -0.144689 noff = 4
+ voffcv = 0 acde = 0.401 moin = 15.773
+ cgsl = {9.82591E-12/sw_func_tox_hv_ratio} cgdl = {9.82591E-12/sw_func_tox_hv_ratio} ijthsrev = 0.1
+ ijthsfwd = 0.1 xjbvs = 1 bvs = 12.69
+ jss = 2.1483E-5 jsws = 4.02E-12 cjs = {sw_psd_nw_cj}
+ mjs = 0.33956 mjsws = 0.24676 cjsws = {9.960545E-11*sw_func_psd_nw_cj}
+ cjswgs = {1.47314E-10*sw_func_psd_nw_cj} mjswgs = 0.81 pbs = 0.6587
+ pbsws = 1 pbswgs = 3 xrcrg1 = 12
+ xrcrg2 = 1 rbpb = 50 rbpd = 50
+ rbps = 50 rbdb = 50 rbsb = 50
+ gbmin = 1E-12 tnom = 30 ute = -1.343412
+ lute = -9.673283E-8 kt1 = -0.569245 lkt1 = -3.613085E-8
+ wkt1 = -5.841868E-8 pkt1 = 2.738055E-14 kt1l = 0
+ kt2 = -0.019032 ua1 = 5.524E-10 ub1 = -3.5909E-18
+ uc1 = -1.092E-10 at = -3.744202E4 lat = 6.13217E-2
+ wat = 0.100378 pat = -9.126851E-8 prt = 0
+ njs = 1.3632 xtis = 10 tpb = 1.671E-3
+ tpbsw = 0 tpbswg = 0 tcj = 9.6E-4
+ tcjsw = 3E-5 tcjswg = 0 tvoff = 0
+ tvfbsdoff = 0 saref = 2.81E-6 sbref = 2.81E-6
+ wlod = 0 ku0 = 7E-8 kvsat = 0.4
+ kvth0 = 3.5E-8 tku0 = 0 llodku0 = 0
+ wlodku0 = 1 llodvth = 0 wlodvth = 1
+ lku0 = 0 wku0 = 0 pku0 = 0
+ lkvth0 = 0 wkvth0 = 6.5E-7 pkvth0 = 0
+ stk2 = 0 lodk2 = 1 steta0 = 0
+ lodeta0 = 1

.model phv_model.41 pmos
+ level = 54 lmin = 6E-7 lmax = 8E-7 wmin = 7.5E-7
+ wmax = 1E-6 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 1.175E-8
+ toxm = 1.175E-8 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 1E23 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {1.2277E-8+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {4.5375E-8-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = -4.7338E-9 dwb = 0 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = -1.17417 lvth0 = 1.495041E-7
+ wvth0 = 2.343035E-7 pvth0 = -1.369277E-13 k1 = -7.79092E-2
+ lk1 = 4.997005E-7 wk1 = 5.136344E-7 pk1 = -3.986646E-13
+ k2 = 0.247926 lk2 = -1.632017E-7 wk2 = -1.885855E-7
+ pk2 = 1.441125E-13 k3 = -2.2405 k3b = -0.172
+ w0 = 0 lpe0 = 0 lpeb = 0
+ vbm = -3 dvtp0 = 0 dvtp1 = 0
+ dvt0 = 4.657 dvt1 = 0.34864 dvt2 = -0.030206
+ dvt0w = -2.2 dvt1w = 1.0163E6 dvt2w = 0
+ vfbsdoff = 0 u0 = 2.10098E-2 lu0 = -5.104018E-9
+ wu0 = -2.349751E-9 pu0 = 3.088513E-15 ua = 1.010545E-10
+ lua = -4.319758E-16 wua = 1.698322E-15 pua = 1.028727E-22
+ ub = 6.222966E-18 lub = -1.619632E-24 wub = -5.304332E-24
+ pub = 1.610198E-30 uc = -7.606797E-12 luc = 5.921598E-18
+ wuc = 7.722576E-18 puc = -7.298289E-24 ud = 0
+ up = 0 lp = 1 eu = 1.67
+ vsat = -9.996654E4 lvsat = 7.90464E-2 wvsat = 0.116426
+ pvsat = -5.119663E-8 a0 = 0.082885 la0 = 6.224159E-7
+ wa0 = 5.813634E-7 pa0 = -5.261002E-13 ags = 5.86162
+ lags = -3.011285E-6 wags = -4.966406E-6 pags = 2.913503E-12
+ b0 = 0 b1 = 0 keta = -0.400154
+ lketa = 1.72131E-7 wketa = 2.946793E-7 pketa = -1.447696E-13
+ a1 = 0 a2 = 0.5 rdsw = 788.47
+ rdswmin = 0 rdw = 0 rdwmin = 0
+ rsw = 0 rswmin = 0 prwb = 0.053538
+ prwg = 0 wr = 1 voff = -0.316616
+ lvoff = 1.490359E-7 wvoff = 2.182203E-7 pvoff = -1.389513E-13
+ voffl = 0 minv = 0 nfactor = 0.822037
+ lnfactor = 2.202105E-7 wnfactor = 4.637291E-7 pnfactor = -2.09428E-14
+ eta0 = 4.90944E-2 leta0 = -9.025504E-8 weta0 = -6.868697E-8
+ peta0 = 1.075111E-13 etab = -4.42921E-2 letab = 2.901684E-8
+ wetab = 2.904094E-8 petab = -2.109155E-14 dsub = -0.289755
+ ldsub = 2.891582E-7 wdsub = 5.249079E-7 pdsub = -2.704077E-13
+ cit = 1E-5 cdsc = 0 cdscb = 0
+ cdscd = 0 pclm = 0.652818 lpclm = 3.173202E-7
+ wpclm = 6.187519E-7 ppclm = -4.025556E-13 pdiblc1 = -1.967614
+ lpdiblc1 = 1.52728E-6 wpdiblc1 = 2.500326E-6 ppdiblc1 = -1.587686E-12
+ pdiblc2 = 1.98826E-2 lpdiblc2 = -6.640821E-12 wpdiblc2 = -1.604376E-8
+ ppdiblc2 = 2.198635E-15 pdiblcb = -0.025 drout = 4.181701
+ ldrout = -2.331051E-6 wdrout = -3.78524E-6 pdrout = 2.443259E-12
+ pscbe1 = 1.834778E9 lpscbe1 = -852.819465 wpscbe1 = -1.354361E3
+ ppscbe1 = 7.783282E-4 pscbe2 = 9.41615E-10 lpscbe2 = 6.776915E-15
+ wpscbe2 = 9.425885E-15 ppscbe2 = -4.618313E-21 pvag = 0
+ delta = 0.01 fprout = 0 pdits = 0
+ pditsl = 0 pditsd = 0 lambda = 0
+ vtl = 0 lc = 5E-9 xn = 3
+ alpha0 = 2.980659E-4 lalpha0 = -1.215876E-10 walpha0 = -2.521328E-10
+ palpha0 = 1.136688E-16 alpha1 = -1.029045E-9 lalpha1 = 5.240412E-16
+ walpha1 = 1.003778E-15 palpha1 = -5.111739E-22 beta0 = 491.501818
+ lbeta0 = -2.234683E-4 wbeta0 = -4.349578E-4 pbeta0 = 2.192627E-10
+ aigbacc = 0.43 bigbacc = 0.054 cigbacc = 0.075
+ nigbacc = 1 aigbinv = 0.35 bigbinv = 0.03
+ cigbinv = 6E-3 eigbinv = 1.1 nigbinv = 3
+ aigc = 0.43 bigc = 0.054 cigc = 0.075
+ aigsd = 0.43 bigsd = 0.054 cigsd = 0.075
+ dlcig = 0 nigc = 1 poxedge = 1
+ pigcd = 1 ntox = 1 toxref = 1.175E-8
+ agidl = -1.168007E-7 lagidl = 1.038082E-13 wagidl = 2.402407E-14
+ pagidl = -3.212626E-20 bgidl = 1.196026E10 lbgidl = -5.649892E3
+ wbgidl = -9.326302E3 pbgidl = 5.088737E-3 cgidl = -6.563258E3
+ lcgidl = 4.020469E-3 wcgidl = 5.767001E-3 pcgidl = -3.118468E-9
+ egidl = -12.304737 legidl = 7.303576E-6 wegidl = 9.55014E-6
+ pegidl = -5.272673E-12 noia = 3E40 noib = 8.53E24
+ noic = 8.4E7 em = 4.1E7 af = 1
+ ef = 0.88 kf = 0 lintnoi = 0
+ tnoia = 1.5 tnoib = 3.5 ntnoi = 1
+ rnoia = 0.577 rnoib = 0.37 xpart = 0
+ cgso = {1.94171E-10/sw_func_tox_hv_ratio} cgdo = {1.94171E-10/sw_func_tox_hv_ratio} cgbo = {0/sw_func_tox_hv_ratio}
+ ckappas = 0.6 cf = 1.2E-11 clc = 1E-7
+ cle = 0.6 dlc = 4.4983E-8 dwc = 0
+ vfbcv = -0.144689 noff = 4 voffcv = 0
+ acde = 0.401 moin = 15.773 cgsl = {9.82591E-12/sw_func_tox_hv_ratio}
+ cgdl = {9.82591E-12/sw_func_tox_hv_ratio} ijthsrev = 0.1 ijthsfwd = 0.1
+ xjbvs = 1 bvs = 12.69 jss = 2.1483E-5
+ jsws = 4.02E-12 cjs = {sw_psd_nw_cj} mjs = 0.33956
+ mjsws = 0.24676 cjsws = {9.960545E-11*sw_func_psd_nw_cj} cjswgs = {1.47314E-10*sw_func_psd_nw_cj}
+ mjswgs = 0.81 pbs = 0.6587 pbsws = 1
+ pbswgs = 3 xrcrg1 = 12 xrcrg2 = 1
+ rbpb = 50 rbpd = 50 rbps = 50
+ rbdb = 50 rbsb = 50 gbmin = 1E-12
+ tnom = 30 ute = -2.042548 lute = 3.991293E-7
+ wute = 2.046858E-7 pute = -1.451734E-13 kt1 = -0.498473
+ lkt1 = -8.632589E-8 wkt1 = -1.063007E-7 pkt1 = 6.134087E-14
+ kt1l = 0 kt2 = -0.019032 ua1 = 5.524E-10
+ ub1 = -1.394971E-17 lub1 = 7.346989E-24 wub1 = 5.829221E-24
+ pub1 = -4.134375E-30 uc1 = -1.092E-10 at = 1.114237E5
+ lat = -4.42613E-2 wat = -6.43416E-2 pat = 2.55587E-8
+ prt = 0 njs = 1.3632 xtis = 10
+ tpb = 1.671E-3 tpbsw = 0 tpbswg = 0
+ tcj = 9.6E-4 tcjsw = 3E-5 tcjswg = 0
+ tvoff = 0 tvfbsdoff = 0 saref = 2.41E-6
+ sbref = 2.41E-6 wlod = 0 ku0 = 7E-8
+ kvsat = 0.4 kvth0 = 3.5E-8 tku0 = 0
+ llodku0 = 0 wlodku0 = 1 llodvth = 0
+ wlodvth = 1 lku0 = 0 wku0 = 0
+ pku0 = 0 lkvth0 = 0 wkvth0 = 6.5E-7
+ pkvth0 = 0 stk2 = 0 lodk2 = 1
+ steta0 = 0 lodeta0 = 1

.model phv_model.42 pmos
+ level = 54 lmin = 5E-7 lmax = 6E-7 wmin = 7.5E-7
+ wmax = 1E-6 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 1.175E-8
+ toxm = 1.175E-8 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 1E23 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {1.2277E-8+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {4.5375E-8-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = -4.7338E-9 dwb = 0 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = -0.369864 lvth0 = -2.600885E-7
+ wvth0 = -4.050835E-7 pvth0 = 1.886802E-13 k1 = 1.98725
+ lk1 = -5.519818E-7 wk1 = -1.055531E-6 pk1 = 4.00433E-13
+ k2 = -0.432333 lk2 = 1.8322E-7 wk2 = 3.55408E-7
+ pk2 = -1.329162E-13 k3 = -2.2405 k3b = -0.172
+ w0 = 0 lpe0 = 0 lpeb = 0
+ vbm = -3 dvtp0 = 0 dvtp1 = 0
+ dvt0 = 4.657 dvt1 = 0.34864 dvt2 = -0.030206
+ dvt0w = -2.2 dvt1w = 1.0163E6 dvt2w = 0
+ vfbsdoff = 0 u0 = -2.783479E-3 lu0 = 7.012723E-9
+ wu0 = 1.370497E-8 pu0 = -5.087352E-15 ua = -2.059636E-9
+ lua = 6.683558E-16 wua = 2.852429E-15 pua = -4.848561E-22
+ ub = -1.478334E-18 lub = 2.302255E-24 wub = 1.13722E-24
+ pub = -1.670162E-30 uc = 5.504698E-11 luc = -2.598484E-17
+ wuc = -4.362526E-17 puc = 1.88506E-23 ud = 0
+ up = 0 lp = 1 eu = 1.67
+ vsat = -6.370146E5 lvsat = 0.352538 wvsat = 0.518097
+ pvsat = -2.557474E-7 a0 = 3.241551 la0 = -9.861349E-7
+ wa0 = -1.856512E-6 pa0 = 7.153876E-13 ags = 9.631748
+ lags = -4.931223E-6 wags = -6.269956E-6 pags = 3.577336E-12
+ b0 = 0 b1 = 0 keta = -0.748699
+ lketa = 3.496278E-7 wketa = 5.084575E-7 pketa = -2.536361E-13
+ a1 = 0 a2 = 0.5 rdsw = 788.47
+ rdswmin = 0 rdw = 0 rdwmin = 0
+ rsw = 0 rswmin = 0 prwb = 0.053538
+ prwg = 0 wr = 1 voff = 0.506417
+ lvoff = -2.700936E-7 wvoff = -4.393931E-7 pvoff = 1.959383E-13
+ voffl = 0 minv = 0 nfactor = 2.445355
+ lnfactor = -6.064644E-7 wnfactor = -4.413273E-7 pnfactor = 4.399572E-13
+ eta0 = -2.340542 leta0 = 1.126667E-6 weta0 = 1.74741E-6
+ peta0 = -8.173364E-13 etab = 0.187474 letab = -8.900992E-8
+ wetab = -1.39174E-7 petab = 6.457189E-14 dsub = 0.176177
+ ldsub = 5.188247E-8 wdsub = 6.782443E-8 pdsub = -3.763793E-14
+ cit = 8.984026E-5 lcit = -4.065865E-11 wcit = -5.791979E-11
+ pcit = 2.949565E-17 cdsc = 0 cdscb = 0
+ cdscd = 0 pclm = 8.606855 lpclm = -3.733273E-6
+ wpclm = -5.489925E-6 ppclm = 2.708288E-12 pdiblc1 = 5.274823
+ lpdiblc1 = -2.160931E-6 wpdiblc1 = -3.695696E-6 ppdiblc1 = 1.567638E-12
+ pdiblc2 = 0.112005 lpdiblc2 = -4.692E-8 wpdiblc2 = -7.856569E-8
+ ppdiblc2 = 3.403792E-14 pdiblcb = 3.16861 lpdiblcb = -1.626346E-6
+ wpdiblcb = -2.316792E-6 ppdiblcb = 1.179826E-12 drout = -6.107704
+ ldrout = 2.908828E-6 wdrout = 5.156255E-6 pdrout = -2.110198E-12
+ pscbe1 = -7.208808E9 lpscbe1 = 3.752627E3 wpscbe1 = 5.519779E3
+ ppscbe1 = -2.722328E-3 pscbe2 = 1.568215E-7 lpscbe2 = -7.26049E-14
+ wpscbe2 = -1.030714E-13 ppscbe2 = 5.267093E-20 pvag = 0
+ delta = 0.01 fprout = 0 pdits = 0
+ pditsl = 0 pditsd = 0 lambda = 0
+ vtl = 0 lc = 5E-9 xn = 3
+ alpha0 = 4.689674E-4 lalpha0 = -2.086192E-10 walpha0 = -3.261105E-10
+ palpha0 = 1.513419E-16 alpha1 = 0 beta0 = 213.737822
+ lbeta0 = -8.201695E-5 wbeta0 = -1.212339E-4 pbeta0 = 5.949887E-11
+ aigbacc = 0.43 bigbacc = 0.054 cigbacc = 0.075
+ nigbacc = 1 aigbinv = 0.35 bigbinv = 0.03
+ cigbinv = 6E-3 eigbinv = 1.1 nigbinv = 3
+ aigc = 0.43 bigc = 0.054 cigc = 0.075
+ aigsd = 0.43 bigsd = 0.054 cigsd = 0.075
+ dlcig = 0 nigc = 1 poxedge = 1
+ pigcd = 1 ntox = 1 toxref = 1.175E-8
+ agidl = 6.395392E-7 lagidl = -2.813579E-13 wagidl = -4.398663E-13
+ pagidl = 2.041099E-19 bgidl = -7.078385E9 lbgidl = 4.045536E3
+ wbgidl = 6.429327E3 pbgidl = -2.934818E-3 cgidl = 1.196635E4
+ lcgidl = -5.415732E-3 wcgidl = -8.071564E-3 pcgidl = 3.928821E-9
+ egidl = 19.250386 legidl = -8.765871E-6 wegidl = -1.329098E-5
+ pegidl = 6.359166E-12 noia = 3E40 noib = 8.53E24
+ noic = 8.4E7 em = 4.1E7 af = 1
+ ef = 0.88 kf = 0 lintnoi = 0
+ tnoia = 1.5 tnoib = 3.5 ntnoi = 1
+ rnoia = 0.577 rnoib = 0.37 xpart = 0
+ cgso = {1.94171E-10/sw_func_tox_hv_ratio} cgdo = {1.94171E-10/sw_func_tox_hv_ratio} cgbo = {0/sw_func_tox_hv_ratio}
+ ckappas = 0.6 cf = 1.2E-11 clc = 1E-7
+ cle = 0.6 dlc = 4.4983E-8 dwc = 0
+ vfbcv = -0.144689 noff = 4 voffcv = 0
+ acde = 0.401 moin = 15.773 cgsl = {9.82591E-12/sw_func_tox_hv_ratio}
+ cgdl = {9.82591E-12/sw_func_tox_hv_ratio} ijthsrev = 0.1 ijthsfwd = 0.1
+ xjbvs = 1 bvs = 12.69 jss = 2.1483E-5
+ jsws = 4.02E-12 cjs = {sw_psd_nw_cj} mjs = 0.33956
+ mjsws = 0.24676 cjsws = {9.960545E-11*sw_func_psd_nw_cj} cjswgs = {1.47314E-10*sw_func_psd_nw_cj}
+ mjswgs = 0.81 pbs = 0.6587 pbsws = 1
+ pbswgs = 3 xrcrg1 = 12 xrcrg2 = 1
+ rbpb = 50 rbpd = 50 rbps = 50
+ rbdb = 50 rbsb = 50 gbmin = 1E-12
+ tnom = 30 ute = -3.181343 lute = 9.790603E-7
+ wute = 1.314321E-6 pute = -7.102554E-13 kt1 = -1.466391
+ lkt1 = 4.065865E-7 wkt1 = 5.933506E-7 pkt1 = -2.949565E-13
+ kt1l = 0 kt2 = -0.019032 ua1 = 5.52E-10
+ ub1 = 5.114485E-18 lub1 = -2.361454E-24 wub1 = -5.653317E-24
+ pub1 = 1.713108E-30 uc1 = -1.092E-10 at = 1.682214E5
+ lat = -7.31856E-2 wat = -0.118408 pat = 5.309218E-8
+ prt = 0 njs = 1.3632 xtis = 10
+ tpb = 1.671E-3 tpbsw = 0 tpbswg = 0
+ tcj = 9.6E-4 tcjsw = 3E-5 tcjswg = 0
+ tvoff = 0 tvfbsdoff = 0 saref = 1.81E-6
+ sbref = 1.81E-6 wlod = 0 ku0 = 7E-8
+ kvsat = 0.4 kvth0 = 3.5E-8 tku0 = 0
+ llodku0 = 0 wlodku0 = 1 llodvth = 0
+ wlodvth = 1 lku0 = 0 wku0 = 0
+ pku0 = 0 lkvth0 = 0 wkvth0 = 6.5E-7
+ pkvth0 = 0 stk2 = 0 lodk2 = 1
+ steta0 = 0 lodeta0 = 1

.model phv_model.43 pmos
+ level = 54 lmin = 8E-6 lmax = 2.02E-5 wmin = 4.2E-7
+ wmax = 7.5E-7 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 1.175E-8
+ toxm = 1.175E-8 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 1E23 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {1.2277E-8+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {4.5375E-8-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = -4.7338E-9 dwb = 0 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = -0.938436 wvth0 = -1.578089E-8
+ k1 = 0.620224 wk1 = -2.566225E-8 k2 = 1.43736E-2
+ wk2 = 7.875275E-9 k3 = -2.2405 k3b = -0.172
+ w0 = 0 lpe0 = 0 lpeb = 0
+ vbm = -3 dvtp0 = 0 dvtp1 = 0
+ dvt0 = 4.657 dvt1 = 0.34864 dvt2 = -0.030206
+ dvt0w = -2.2 dvt1w = 1.0163E6 dvt2w = 0
+ vfbsdoff = 0 u0 = 1.65676E-2 wu0 = 1.476318E-9
+ ua = 2.294564E-9 wua = -3.198171E-17 ub = 1.992005E-19
+ wub = 3.51352E-26 uc = -6.136091E-11 wuc = 1.179019E-17
+ ud = 0 up = 0 lp = 1
+ eu = 1.67 vsat = 8.0156E4 a0 = 0.938091
+ wa0 = -2.297201E-8 ags = 0.159749 wags = -1.607053E-8
+ b0 = -7.217489E-9 wb0 = 5.235898E-15 b1 = -5.397359E-10
+ wb1 = 3.915492E-16 keta = -1.18117E-2 wketa = 2.633249E-9
+ a1 = 0 a2 = 0.5 rdsw = 788.47
+ rdswmin = 0 rdw = 0 rdwmin = 0
+ rsw = 0 rswmin = 0 prwb = 0.053538
+ prwg = 0 wr = 1 voff = -8.43405E-2
+ wvoff = -1.693161E-8 voffl = 0 minv = 0
+ nfactor = 1.470232 wnfactor = 9.313866E-8 eta0 = 0.08
+ etab = -0.07 dsub = 0.56 cit = 7.995803E-6
+ wcit = -2.173293E-12 cdsc = 0 cdscb = 0
+ cdscd = 0 pclm = 0.083531 pdiblc1 = 0.39
+ pdiblc2 = 7.967041E-4 wpdiblc2 = 1.916166E-9 pdiblcb = -0.025
+ drout = 0.56 pscbe1 = 2.243792E8 wpscbe1 = 0.245487
+ pscbe2 = 1.5E-8 pvag = 0 delta = 0.01
+ fprout = 0 pdits = 0 pditsl = 0
+ pditsd = 0 lambda = 0 vtl = 0
+ lc = 5E-9 xn = 3 alpha0 = 1.412258E-4
+ walpha0 = -5.584715E-11 alpha1 = -1.198321E-10 walpha1 = 8.693173E-17
+ beta0 = 82.226349 wbeta0 = -3.132974E-5 aigbacc = 0.43
+ bigbacc = 0.054 cigbacc = 0.075 nigbacc = 1
+ aigbinv = 0.35 bigbinv = 0.03 cigbinv = 6E-3
+ eigbinv = 1.1 nigbinv = 3 aigc = 0.43
+ bigc = 0.054 cigc = 0.075 aigsd = 0.43
+ bigsd = 0.054 cigsd = 0.075 dlcig = 0
+ nigc = 1 poxedge = 1 pigcd = 1
+ ntox = 1 toxref = 1.175E-8 agidl = -3.991606E-8
+ wagidl = 4.346587E-14 bgidl = 1.78451E9 wbgidl = -191.59754
+ cgidl = 1.298143E3 wcgidl = 7.389197E-5 egidl = 0.944663
+ wegidl = 4.173287E-7 noia = 3E40 noib = 8.53E24
+ noic = 8.4E7 em = 4.1E7 af = 1
+ ef = 0.88 kf = 0 lintnoi = 0
+ tnoia = 1.5 tnoib = 3.5 ntnoi = 1
+ rnoia = 0.577 rnoib = 0.37 xpart = 0
+ cgso = {1.94171E-10/sw_func_tox_hv_ratio} cgdo = {1.94171E-10/sw_func_tox_hv_ratio} cgbo = {0/sw_func_tox_hv_ratio}
+ ckappas = 0.6 cf = 1.2E-11 clc = 1E-7
+ cle = 0.6 dlc = 4.4983E-8 dwc = 0
+ vfbcv = -0.144689 noff = 4 voffcv = 0
+ acde = 0.401 moin = 15.773 cgsl = {9.82591E-12/sw_func_tox_hv_ratio}
+ cgdl = {9.82591E-12/sw_func_tox_hv_ratio} ijthsrev = 0.1 ijthsfwd = 0.1
+ xjbvs = 1 bvs = 12.69 jss = 2.1483E-5
+ jsws = 4.02E-12 cjs = {sw_psd_nw_cj} mjs = 0.33956
+ mjsws = 0.24676 cjsws = {9.960545E-11*sw_func_psd_nw_cj} cjswgs = {1.47314E-10*sw_func_psd_nw_cj}
+ mjswgs = 0.81 pbs = 0.6587 pbsws = 1
+ pbswgs = 3 xrcrg1 = 12 xrcrg2 = 1
+ rbpb = 50 rbpd = 50 rbps = 50
+ rbdb = 50 rbsb = 50 gbmin = 1E-12
+ tnom = 30 ute = -1.5561 kt1 = -0.567983
+ wkt1 = 8.693173E-9 kt1l = 0 kt2 = -0.019032
+ ua1 = 2.2096E-11 ub1 = -3.0767E-18 uc1 = -1.092E-10
+ at = 1.5109E5 prt = 0 njs = 1.3632
+ xtis = 10 tpb = 1.671E-3 tpbsw = 0
+ tpbswg = 0 tcj = 9.6E-4 tcjsw = 3E-5
+ tcjswg = 0 tvoff = 0 tvfbsdoff = 0
+ saref = 3E-6 sbref = 3E-6 wlod = 0
+ ku0 = 7E-8 kvsat = 0.4 kvth0 = 3.5E-8
+ tku0 = 0 llodku0 = 0 wlodku0 = 1
+ llodvth = 0 wlodvth = 1 lku0 = 0
+ wku0 = 0 pku0 = 0 lkvth0 = 0
+ wkvth0 = 6.5E-7 pkvth0 = 0 stk2 = 0
+ lodk2 = 1 steta0 = 0 lodeta0 = 1

.model phv_model.44 pmos
+ level = 54 lmin = 4E-6 lmax = 8E-6 wmin = 4.2E-7
+ wmax = 7.5E-7 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 1.175E-8
+ toxm = 1.175E-8 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 1E23 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {1.2277E-8+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {4.5375E-8-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = -4.7338E-9 dwb = 0 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = -0.971394 lvth0 = 2.606723E-7
+ wvth0 = -1.827318E-9 pvth0 = -1.103623E-13 k1 = 0.617872
+ lk1 = 1.860563E-8 wk1 = -3.831271E-8 pk1 = 1.000557E-13
+ k2 = 1.24447E-2 lk2 = 1.525567E-8 wk2 = 1.378171E-8
+ pk2 = -4.671545E-14 k3 = -2.2405 k3b = -0.172
+ w0 = 0 lpe0 = 0 lpeb = 0
+ vbm = -3 dvtp0 = 0 dvtp1 = 0
+ dvt0 = 4.657 dvt1 = 0.34864 dvt2 = -0.030206
+ dvt0w = -2.2 dvt1w = 1.0163E6 dvt2w = 0
+ vfbsdoff = 0 u0 = 1.88178E-2 lu0 = -1.779772E-8
+ wu0 = 3.784804E-10 pu0 = 8.683073E-15 ua = 2.78929E-9
+ lua = -3.91291E-15 wua = -1.896852E-16 pua = 1.247317E-21
+ ub = 2.208971E-19 lub = -1.716041E-25 wub = -7.344432E-26
+ pub = 8.587826E-31 uc = -8.9242E-11 luc = 2.205185E-16
+ wuc = 2.123518E-17 puc = -7.470282E-23 ud = 0
+ up = 0 lp = 1 eu = 1.67
+ vsat = 4.099118E4 lvsat = 0.309764 a0 = 0.93973
+ la0 = -1.296247E-8 wa0 = 3.433091E-9 pa0 = -2.088446E-13
+ ags = 0.153997 lags = 4.549451E-8 wags = -1.214523E-8
+ pags = -3.104616E-14 b0 = 9.710824E-10 lb0 = -6.476546E-14
+ wb0 = -7.044678E-16 pb0 = 4.698384E-20 b1 = 6.7515E-9
+ lb1 = -5.766821E-14 wb1 = -4.897849E-15 pb1 = 4.183517E-20
+ keta = -8.16798E-3 lketa = -2.881937E-8 wketa = 1.156399E-9
+ pketa = 1.168078E-14 a1 = 0 a2 = 0.5
+ rdsw = 788.47 rdswmin = 0 rdw = 0
+ rdwmin = 0 rsw = 0 rswmin = 0
+ prwb = 0.053538 prwg = 0 wr = 1
+ voff = -0.129461 lvoff = 3.568667E-7 wvoff = 8.278535E-9
+ pvoff = -1.993933E-13 voffl = 0 minv = 0
+ nfactor = 0.817604 lnfactor = 5.1618E-6 wnfactor = 5.230676E-7
+ pnfactor = -3.400415E-12 eta0 = 0.08 etab = -0.07
+ dsub = 0.56 cit = 1.814048E-7 lcit = 6.180603E-11
+ wcit = -4.930659E-14 pcit = -1.679914E-17 cdsc = 0
+ cdscb = 0 cdscd = 0 pclm = -0.279769
+ lpclm = 2.873436E-6 wpclm = -3.249694E-7 ppclm = 2.570263E-12
+ pdiblc1 = 0.39 pdiblc2 = 3.145998E-4 lpdiblc2 = 3.813083E-9
+ wpdiblc2 = 3.788859E-9 ppdiblc2 = -1.48116E-14 pdiblcb = -0.025
+ drout = 0.56 pscbe1 = 2.236482E8 lpscbe1 = 5.782159
+ wpscbe1 = 0.534026 ppscbe1 = -2.28213E-6 pscbe2 = 1.5E-8
+ pvag = 0 delta = 0.01 fprout = 0
+ pdits = 0 pditsl = 0 pditsd = 0
+ lambda = 0 vtl = 0 lc = 5E-9
+ xn = 3 alpha0 = 3.050831E-4 lalpha0 = -1.295988E-9
+ walpha0 = -1.291696E-10 palpha0 = 5.799253E-16 alpha1 = -4.517902E-10
+ lalpha1 = 2.62554E-15 walpha1 = 2.568507E-16 palpha1 = -1.343931E-21
+ beta0 = 199.431203 lbeta0 = -9.270025E-4 wbeta0 = -9.0804E-5
+ pbeta0 = 4.703968E-10 aigbacc = 0.43 bigbacc = 0.054
+ cigbacc = 0.075 nigbacc = 1 aigbinv = 0.35
+ bigbinv = 0.03 cigbinv = 6E-3 eigbinv = 1.1
+ nigbinv = 3 aigc = 0.43 bigc = 0.054
+ cigc = 0.075 aigsd = 0.43 bigsd = 0.054
+ cigsd = 0.075 dlcig = 0 nigc = 1
+ poxedge = 1 pigcd = 1 ntox = 1
+ toxref = 1.175E-8 agidl = -7.651308E-8 lagidl = 2.89455E-13
+ wagidl = 6.03728E-14 pagidl = -1.337212E-19 bgidl = 2.22284E9
+ lbgidl = -3.466861E3 wbgidl = -475.479921 pbgidl = 2.245297E-3
+ cgidl = 2.915159E3 lcgidl = -1.27894E-2 wcgidl = -4.554055E-4
+ pcgidl = 4.186346E-9 egidl = -0.872368 legidl = 1.437136E-5
+ wegidl = 1.395127E-6 pegidl = -7.733652E-12 noia = 3E40
+ noib = 8.53E24 noic = 8.4E7 em = 4.1E7
+ af = 1 ef = 0.88 kf = 0
+ lintnoi = 0 tnoia = 1.5 tnoib = 3.5
+ ntnoi = 1 rnoia = 0.577 rnoib = 0.37
+ xpart = 0 cgso = {1.94171E-10/sw_func_tox_hv_ratio} cgdo = {1.94171E-10/sw_func_tox_hv_ratio}
+ cgbo = {0/sw_func_tox_hv_ratio} ckappas = 0.6 cf = 1.2E-11
+ clc = 1E-7 cle = 0.6 dlc = 4.4983E-8
+ dwc = 0 vfbcv = -0.144689 noff = 4
+ voffcv = 0 acde = 0.401 moin = 15.773
+ cgsl = {9.82591E-12/sw_func_tox_hv_ratio} cgdl = {9.82591E-12/sw_func_tox_hv_ratio} ijthsrev = 0.1
+ ijthsfwd = 0.1 xjbvs = 1 bvs = 12.69
+ jss = 2.1483E-5 jsws = 4.02E-12 cjs = {sw_psd_nw_cj}
+ mjs = 0.33956 mjsws = 0.24676 cjsws = {9.960545E-11*sw_func_psd_nw_cj}
+ cjswgs = {1.47314E-10*sw_func_psd_nw_cj} mjswgs = 0.81 pbs = 0.6587
+ pbsws = 1 pbswgs = 3 xrcrg1 = 12
+ xrcrg2 = 1 rbpb = 50 rbpd = 50
+ rbps = 50 rbdb = 50 rbsb = 50
+ gbmin = 1E-12 tnom = 30 ute = -1.735971
+ lute = 1.422643E-6 wute = 2.718703E-8 pute = -2.15029E-13
+ kt1 = -0.548437 lkt1 = -1.545962E-7 wkt1 = 8.693173E-9
+ kt1l = 0 kt2 = -0.019032 ua1 = 2.2096E-11
+ ub1 = -3.738243E-18 lub1 = 5.232308E-24 uc1 = -1.092E-10
+ at = 8.408545E4 lat = 0.529956 prt = 0
+ njs = 1.3632 xtis = 10 tpb = 1.671E-3
+ tpbsw = 0 tpbswg = 0 tcj = 9.6E-4
+ tcjsw = 3E-5 tcjswg = 0 tvoff = 0
+ tvfbsdoff = 0 saref = 3E-6 sbref = 3E-6
+ wlod = 0 ku0 = 7E-8 kvsat = 0.4
+ kvth0 = 3.5E-8 tku0 = 0 llodku0 = 0
+ wlodku0 = 1 llodvth = 0 wlodvth = 1
+ lku0 = 0 wku0 = 0 pku0 = 0
+ lkvth0 = 0 wkvth0 = 6.5E-7 pkvth0 = 0
+ stk2 = 0 lodk2 = 1 steta0 = 0
+ lodeta0 = 1

.model phv_model.45 pmos
+ level = 54 lmin = 2E-6 lmax = 4E-6 wmin = 4.2E-7
+ wmax = 7.5E-7 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 1.175E-8
+ toxm = 1.175E-8 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 1E23 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {1.2277E-8+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {4.5375E-8-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = -4.7338E-9 dwb = 0 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = -0.957508 lvth0 = 2.063898E-7
+ wvth0 = -9.836063E-9 pvth0 = -7.905411E-14 k1 = 0.718665
+ lk1 = -3.754202E-7 wk1 = -5.10416E-8 pk1 = 1.498161E-13
+ k2 = -1.94046E-2 lk2 = 1.397629E-7 wk2 = 1.675726E-8
+ pk2 = -5.834761E-14 k3 = -2.2405 k3b = -0.172
+ w0 = 0 lpe0 = 0 lpeb = 0
+ vbm = -3 dvtp0 = 0 dvtp1 = 0
+ dvt0 = 4.657 dvt1 = 0.34864 dvt2 = -0.030206
+ dvt0w = -2.2 dvt1w = 1.0163E6 dvt2w = 0
+ vfbsdoff = 0 u0 = 1.59226E-2 lu0 = -6.479685E-9
+ wu0 = 1.98937E-9 pu0 = 2.385703E-15 ua = 1.473554E-9
+ lua = 1.230631E-15 wua = 3.130331E-16 pua = -7.179348E-22
+ ub = 1.663508E-18 lub = -5.811133E-24 wub = -4.929998E-25
+ pub = 2.49893E-30 uc = -7.14578E-11 luc = 1.509956E-16
+ wuc = 1.137541E-17 puc = -3.615849E-23 ud = 0
+ up = 0 lp = 1 eu = 1.67
+ vsat = 3.045246E5 lvsat = -0.720454 wvsat = -7.68876E-2
+ pvsat = 3.00573E-7 a0 = 1.285454 la0 = -1.364484E-6
+ wa0 = -2.144417E-7 pa0 = 6.428824E-13 ags = -0.46932
+ lags = 2.482198E-6 wags = 2.366052E-7 pags = -1.003474E-12
+ b0 = -1.826671E-7 lb0 = 6.531219E-13 wb0 = 8.631717E-14
+ pb0 = -2.932055E-19 b1 = -8.625444E-9 lb1 = 2.444108E-15
+ wb1 = 5.987138E-15 pb1 = -7.169632E-22 keta = 3.73733E-2
+ lketa = -2.068515E-7 wketa = -1.529255E-8 pketa = 7.598382E-14
+ a1 = 0 a2 = 0.5 rdsw = 788.47
+ rdswmin = 0 rdw = 0 rdwmin = 0
+ rsw = 0 rswmin = 0 prwb = 0.053538
+ prwg = 0 wr = 1 voff = -7.91136E-2
+ lvoff = 1.600473E-7 wvoff = -2.780278E-8 pvoff = -5.834242E-14
+ voffl = 0 minv = 0 nfactor = 1.770907
+ lnfactor = 1.435099E-6 wnfactor = -2.164559E-7 pnfactor = -5.094332E-13
+ eta0 = 0.59099 leta0 = -1.997587E-6 weta0 = -3.56845E-7
+ peta0 = 1.394996E-12 etab = -1.345404 letab = 4.985874E-6
+ wetab = 8.767598E-7 petab = -3.427473E-12 dsub = 0.72896
+ ldsub = -6.605084E-7 wdsub = 4.643608E-8 pdsub = -1.815302E-13
+ cit = 1.599161E-5 wcit = -4.346587E-12 cdsc = 0
+ cdscb = 0 cdscd = 0 pclm = 0.575333
+ lpclm = -4.693714E-7 wpclm = 6.733574E-8 ppclm = 1.036644E-12
+ pdiblc1 = 0.282569 lpdiblc1 = 4.199759E-7 wpdiblc1 = -3.052813E-8
+ ppdiblc1 = 1.193421E-13 pdiblc2 = -2.643173E-4 lpdiblc2 = 6.076215E-9
+ wpdiblc2 = 6.146486E-10 ppdiblc2 = -2.402815E-15 pdiblcb = -0.025
+ drout = 0.555877 ldrout = 1.611718E-8 wdrout = 9.589951E-8
+ pdrout = -3.748952E-13 pscbe1 = 1.913435E8 lpscbe1 = 132.069011
+ wpscbe1 = -12.299451 ppscbe1 = 4.788714E-5 pscbe2 = 1.57562E-8
+ lpscbe2 = -2.892729E-15 wpscbe2 = -2.015134E-16 ppscbe2 = 7.626931E-22
+ pvag = 0 delta = 0.01 fprout = 0
+ pdits = 0 pditsl = 0 pditsd = 0
+ lambda = 0 vtl = 0 lc = 5E-9
+ xn = 3 alpha0 = -4.507122E-5 lalpha0 = 7.285291E-11
+ walpha0 = 3.269681E-11 palpha0 = -5.285085E-17 alpha1 = 2.198321E-10
+ walpha1 = -8.693173E-17 beta0 = -39.635919 lbeta0 = 7.570653E-6
+ wbeta0 = 3.093006E-5 pbeta0 = -5.4921E-12 aigbacc = 0.43
+ bigbacc = 0.054 cigbacc = 0.075 nigbacc = 1
+ aigbinv = 0.35 bigbinv = 0.03 cigbinv = 6E-3
+ eigbinv = 1.1 nigbinv = 3 aigc = 0.43
+ bigc = 0.054 cigc = 0.075 aigsd = 0.43
+ bigsd = 0.054 cigsd = 0.075 dlcig = 0
+ nigc = 1 poxedge = 1 pigcd = 1
+ ntox = 1 toxref = 1.175E-8 agidl = 7.34263E-8
+ lagidl = -2.966955E-13 wagidl = -5.695988E-15 pagidl = 1.245582E-19
+ bgidl = 2.247804E9 lbgidl = -3.564453E3 wbgidl = -255.242176
+ pbgidl = 1.384332E-3 cgidl = -2.883439E3 lcgidl = 9.878783E-3
+ wcgidl = 1.6329E-3 pcgidl = -3.977361E-9 egidl = 5.260082
+ legidl = -9.601922E-6 wegidl = -1.609931E-6 pegidl = 4.013871E-12
+ noia = 3E40 noib = 8.53E24 noic = 8.4E7
+ em = 4.1E7 af = 1 ef = 0.88
+ kf = 0 lintnoi = 0 tnoia = 1.5
+ tnoib = 3.5 ntnoi = 1 rnoia = 0.577
+ rnoib = 0.37 xpart = 0 cgso = {1.94171E-10/sw_func_tox_hv_ratio}
+ cgdo = {1.94171E-10/sw_func_tox_hv_ratio} cgbo = {0/sw_func_tox_hv_ratio} ckappas = 0.6
+ cf = 1.2E-11 clc = 1E-7 cle = 0.6
+ dlc = 4.4983E-8 dwc = 0 vfbcv = -0.144689
+ noff = 4 voffcv = 0 acde = 0.401
+ moin = 15.773 cgsl = {9.82591E-12/sw_func_tox_hv_ratio} cgdl = {9.82591E-12/sw_func_tox_hv_ratio}
+ ijthsrev = 0.1 ijthsfwd = 0.1 xjbvs = 1
+ bvs = 12.69 jss = 2.1483E-5 jsws = 4.02E-12
+ cjs = {sw_psd_nw_cj} mjs = 0.33956 mjsws = 0.24676
+ cjsws = {9.960545E-11*sw_func_psd_nw_cj} cjswgs = {1.47314E-10*sw_func_psd_nw_cj} mjswgs = 0.81
+ pbs = 0.6587 pbsws = 1 pbswgs = 3
+ xrcrg1 = 12 xrcrg2 = 1 rbpb = 50
+ rbpd = 50 rbps = 50 rbdb = 50
+ rbsb = 50 gbmin = 1E-12 tnom = 30
+ ute = -1.183669 lute = -7.364421E-7 wute = -1.371953E-7
+ pute = 4.275826E-13 kt1 = -0.462053 lkt1 = -4.922933E-7
+ wkt1 = -3.280043E-8 pkt1 = 1.622089E-13 kt1l = 0
+ kt2 = -0.019032 ua1 = -4.841455E-10 lua1 = 1.979024E-15
+ ub1 = -8.196953E-19 lub1 = -6.177024E-24 wub1 = -3.214094E-25
+ pub1 = 1.25647E-30 uc1 = -1.092E-10 at = 5.667894E5
+ lat = -1.357055 wat = -0.123817 pat = 4.840313E-7
+ prt = 0 njs = 1.3632 xtis = 10
+ tpb = 1.671E-3 tpbsw = 0 tpbswg = 0
+ tcj = 9.6E-4 tcjsw = 3E-5 tcjswg = 0
+ tvoff = 0 tvfbsdoff = 0 saref = 3E-6
+ sbref = 3E-6 wlod = 0 ku0 = 7E-8
+ kvsat = 0.4 kvth0 = 3.5E-8 tku0 = 0
+ llodku0 = 0 wlodku0 = 1 llodvth = 0
+ wlodvth = 1 lku0 = 0 wku0 = 0
+ pku0 = 0 lkvth0 = 0 wkvth0 = 6.5E-7
+ pkvth0 = 0 stk2 = 0 lodk2 = 1
+ steta0 = 0 lodeta0 = 1

.model phv_model.46 pmos
+ level = 54 lmin = 1E-6 lmax = 2E-6 wmin = 4.2E-7
+ wmax = 7.5E-7 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 1.175E-8
+ toxm = 1.175E-8 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 1E23 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {1.2277E-8+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {4.5375E-8-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = -4.7338E-9 dwb = 0 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = -0.832564 lvth0 = -3.215879E-8
+ wvth0 = -7.120163E-8 pvth0 = 3.81081E-14 k1 = 0.51221
+ lk1 = 1.875439E-8 wk1 = 3.455295E-8 pk1 = -1.36053E-14
+ k2 = 5.97119E-2 lk2 = -1.129044E-8 wk2 = -1.83759E-8
+ pk2 = 8.730371E-15 k3 = -2.2405 k3b = -0.172
+ w0 = 0 lpe0 = 0 lpeb = 0
+ vbm = -3 dvtp0 = 0 dvtp1 = 0
+ dvt0 = 4.657 dvt1 = 0.34864 dvt2 = -0.030206
+ dvt0w = -2.2 dvt1w = 1.0163E6 dvt2w = 0
+ vfbsdoff = 0 u0 = 1.02573E-2 lu0 = 4.336748E-9
+ wu0 = 5.017594E-9 pu0 = -3.395934E-15 ua = 1.9017E-9
+ lua = 4.131933E-16 wua = 9.409378E-17 pua = -2.99925E-22
+ ub = -1.959625E-18 lub = 1.106334E-24 wub = 1.21326E-24
+ pub = -7.587472E-31 uc = 1.547479E-11 luc = -1.498043E-17
+ wuc = -1.32552E-17 puc = 1.086749E-23 ud = 0
+ up = 0 lp = 1 eu = 1.67
+ vsat = -1.804256E5 lvsat = 0.205437 wvsat = 0.137937
+ pvsat = -1.095804E-7 a0 = 0.302071 la0 = 5.13041E-7
+ wa0 = 3.172152E-7 pa0 = -3.721835E-13 ags = 0.861414
+ lags = -5.850755E-8 wags = -3.112108E-7 pags = 4.244407E-14
+ b0 = 1.028564E-7 lb0 = 1.079863E-13 wb0 = -4.155235E-14
+ pb0 = -4.907062E-20 b1 = 4.154673E-8 lb1 = -9.334711E-14
+ wb1 = -3.02823E-14 pb1 = 6.853045E-20 keta = -8.40144E-2
+ lketa = 2.490793E-8 wketa = 3.095685E-8 pketa = -1.231784E-14
+ a1 = 0 a2 = 0.5 rdsw = 788.47
+ rdswmin = 0 rdw = 0 rdwmin = 0
+ rsw = 0 rswmin = 0 prwb = 0.053538
+ prwg = 0 wr = 1 voff = 0.054486
+ lvoff = -9.502778E-8 wvoff = -9.446768E-8 pvoff = 6.893753E-14
+ voffl = 0 minv = 0 nfactor = 3.30842
+ lnfactor = -1.500398E-6 wnfactor = -9.730359E-7 pnfactor = 9.350673E-13
+ eta0 = -0.628232 leta0 = 3.302127E-7 weta0 = 5.150328E-7
+ peta0 = -2.696364E-13 etab = 2.424995 letab = -2.212762E-6
+ wetab = -1.75634E-6 petab = 1.599773E-12 dsub = 0.392068
+ ldsub = -1.729668E-8 wdsub = -5.521538E-8 pdsub = 1.254781E-14
+ cit = 1.599161E-5 wcit = -4.346587E-12 cdsc = 0
+ cdscb = 0 cdscd = 0 pclm = -0.651102
+ lpclm = 1.872199E-6 wpclm = 1.321662E-6 ppclm = -1.358179E-12
+ pdiblc1 = 0.325131 lpdiblc1 = 3.387147E-7 wpdiblc1 = 1.606785E-7
+ ppdiblc1 = -2.457192E-13 pdiblc2 = 2.790262E-3 lpdiblc2 = 2.442587E-10
+ wpdiblc2 = -5.510544E-10 ppdiblc2 = -1.771965E-16 pdiblcb = -0.025
+ drout = 1.180624 ldrout = -1.17668E-6 wdrout = -5.475537E-7
+ pdrout = 8.536178E-13 pscbe1 = 2.78102E8 lpscbe1 = -33.574553
+ wpscbe1 = 2.50818E-2 ppscbe1 = 2.435653E-5 pscbe2 = 1.439587E-8
+ lpscbe2 = -2.955188E-16 wpscbe2 = 8.567276E-17 ppscbe2 = 2.143829E-22
+ pvag = 0 delta = 0.01 fprout = 0
+ pdits = 0 pditsl = 0 pditsd = 0
+ lambda = 0 vtl = 0 lc = 5E-9
+ xn = 3 alpha0 = -1.721933E-6 lalpha0 = -9.911722E-12
+ walpha0 = 1.249242E-12 palpha0 = 7.190419E-18 alpha1 = 2.198321E-10
+ walpha1 = -8.693173E-17 beta0 = -30.288326 lbeta0 = -1.027624E-5
+ wbeta0 = 2.414888E-5 pbeta0 = 7.454856E-12 aigbacc = 0.43
+ bigbacc = 0.054 cigbacc = 0.075 nigbacc = 1
+ aigbinv = 0.35 bigbinv = 0.03 cigbinv = 6E-3
+ eigbinv = 1.1 nigbinv = 3 aigc = 0.43
+ bigc = 0.054 cigc = 0.075 aigsd = 0.43
+ bigsd = 0.054 cigsd = 0.075 dlcig = 0
+ nigc = 1 poxedge = 1 pigcd = 1
+ ntox = 1 toxref = 1.175E-8 agidl = -1.022388E-7
+ lagidl = 3.869299E-14 wagidl = 7.424531E-14 pagidl = -2.806968E-20
+ bgidl = 6.161287E8 lbgidl = -449.176321 wbgidl = 299.153086
+ pbgidl = 3.258532E-4 cgidl = 3.4762E3 lcgidl = -2.263358E-3
+ wcgidl = -8.644426E-4 pcgidl = 7.906896E-10 egidl = -0.545256
+ legidl = 1.48192E-6 wegidl = 1.055473E-6 pegidl = -1.075053E-12
+ noia = 3E40 noib = 8.53E24 noic = 8.4E7
+ em = 4.1E7 af = 1 ef = 0.88
+ kf = 0 lintnoi = 0 tnoia = 1.5
+ tnoib = 3.5 ntnoi = 1 rnoia = 0.577
+ rnoib = 0.37 xpart = 0 cgso = {1.94171E-10/sw_func_tox_hv_ratio}
+ cgdo = {1.94171E-10/sw_func_tox_hv_ratio} cgbo = {0/sw_func_tox_hv_ratio} ckappas = 0.6
+ cf = 1.2E-11 clc = 1E-7 cle = 0.6
+ dlc = 4.4983E-8 dwc = 0 vfbcv = -0.144689
+ noff = 4 voffcv = 0 acde = 0.401
+ moin = 15.773 cgsl = {9.82591E-12/sw_func_tox_hv_ratio} cgdl = {9.82591E-12/sw_func_tox_hv_ratio}
+ ijthsrev = 0.1 ijthsfwd = 0.1 xjbvs = 1
+ bvs = 12.69 jss = 2.1483E-5 jsws = 4.02E-12
+ cjs = {sw_psd_nw_cj} mjs = 0.33956 mjsws = 0.24676
+ cjsws = {9.960545E-11*sw_func_psd_nw_cj} cjswgs = {1.47314E-10*sw_func_psd_nw_cj} mjswgs = 0.81
+ pbs = 0.6587 pbsws = 1 pbswgs = 3
+ xrcrg1 = 12 xrcrg2 = 1 rbpb = 50
+ rbpd = 50 rbps = 50 rbdb = 50
+ rbsb = 50 gbmin = 1E-12 tnom = 30
+ ute = -1.678132 lute = 2.076108E-7 wute = 1.656425E-7
+ pute = -1.506104E-13 kt1 = -0.776557 lkt1 = 1.08174E-7
+ wkt1 = 9.326123E-8 pkt1 = -7.847436E-14 kt1l = 0
+ kt2 = -0.019032 ua1 = 5.524E-10 ub1 = -3.719748E-18
+ lub1 = -6.400986E-25 wub1 = 9.347228E-26 pub1 = 4.643569E-31
+ uc1 = -1.092E-10 at = -3.23981E5 lat = 0.343649
+ wat = 0.263442 pat = -2.553435E-7 prt = 0
+ njs = 1.3632 xtis = 10 tpb = 1.671E-3
+ tpbsw = 0 tpbswg = 0 tcj = 9.6E-4
+ tcjsw = 3E-5 tcjswg = 0 tvoff = 0
+ tvfbsdoff = 0 saref = 3E-6 sbref = 3E-6
+ wlod = 0 ku0 = 7E-8 kvsat = 0.4
+ kvth0 = 3.5E-8 tku0 = 0 llodku0 = 0
+ wlodku0 = 1 llodvth = 0 wlodvth = 1
+ lku0 = 0 wku0 = 0 pku0 = 0
+ lkvth0 = 0 wkvth0 = 6.5E-7 pkvth0 = 0
+ stk2 = 0 lodk2 = 1 steta0 = 0
+ lodeta0 = 1

.model phv_model.47 pmos
+ level = 54 lmin = 8E-7 lmax = 1E-6 wmin = 4.2E-7
+ wmax = 7.5E-7 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 1.175E-8
+ toxm = 1.175E-8 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 1E23 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {1.2277E-8+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {4.5375E-8-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = -4.7338E-9 dwb = 0 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = -0.887288 lvth0 = 1.759908E-8
+ wvth0 = -1.983558E-8 pvth0 = -8.596481E-15 k1 = 0.291838
+ lk1 = 2.191277E-7 wk1 = 1.94421E-7 pk1 = -1.589653E-13
+ k2 = 0.10489 lk2 = -5.236829E-8 wk2 = -5.76397E-8
+ pk2 = 4.443098E-14 k3 = -2.2405 k3b = -0.172
+ w0 = 0 lpe0 = 0 lpeb = 0
+ vbm = -3 dvtp0 = 0 dvtp1 = 0
+ dvt0 = 4.657 dvt1 = 0.34864 dvt2 = -0.030206
+ dvt0w = -2.2 dvt1w = 1.0163E6 dvt2w = 0
+ vfbsdoff = 0 u0 = 0.016251 lu0 = -1.113005E-9
+ wu0 = 9.555379E-10 pu0 = 2.974906E-16 ua = 1.513593E-9
+ lua = 7.660799E-16 wua = 3.70649E-16 pua = -5.513829E-22
+ ub = 1.102139E-18 lub = -1.677574E-24 wub = -9.02532E-25
+ pub = 1.165037E-30 uc = -1.253427E-12 luc = 2.297031E-19
+ wuc = -1.119781E-18 puc = -1.666372E-25 ud = 0
+ up = 0 lp = 1 eu = 1.67
+ vsat = -3.375844E4 lvsat = 7.20803E-2 wvsat = 6.73596E-2
+ pvsat = -4.540814E-8 a0 = 1.426853 la0 = -5.096676E-7
+ wa0 = -4.987539E-7 pa0 = 3.697364E-13 ags = 1.977716
+ lags = -1.073505E-6 wags = -1.121028E-6 pags = 7.787699E-13
+ b0 = 1.007542E-6 lb0 = -7.145994E-13 wb0 = -4.342605E-13
+ pb0 = 3.079992E-19 b1 = -2.778537E-7 lb1 = 1.970678E-13
+ wb1 = 2.049814E-13 pb1 = -1.45383E-19 keta = -0.128994
+ lketa = 6.580551E-8 wketa = 6.991258E-8 pketa = -4.773834E-14
+ a1 = 0 a2 = 0.5 rdsw = 788.47
+ rdswmin = 0 rdw = 0 rdwmin = 0
+ rsw = 0 rswmin = 0 prwb = 0.053538
+ prwg = 0 wr = 1 voff = -0.104793
+ lvoff = 4.979679E-8 wvoff = 2.108076E-8 pvoff = -3.612489E-14
+ voffl = 0 minv = 0 nfactor = 1.17715
+ lnfactor = 4.374592E-7 wnfactor = 4.134667E-7 pnfactor = -3.256103E-13
+ eta0 = 0.595726 leta0 = -7.826716E-7 weta0 = -4.059707E-7
+ peta0 = 5.67786E-13 etab = -5.360226E-3 letab = -2.960791E-9
+ wetab = 7.396108E-10 petab = 2.147894E-15 dsub = 1.226708
+ ldsub = -7.761929E-7 wdsub = -6.607015E-7 pdsub = 5.63086E-13
+ cit = 1.599161E-5 wcit = -4.346587E-12 cdsc = 0
+ cdscb = 0 cdscd = 0 pclm = 1.501257
+ lpclm = -8.483355E-8 wpclm = -2.397579E-7 ppclm = 6.154216E-14
+ pdiblc1 = 0.617252 lpdiblc1 = 7.310333E-8 wpdiblc1 = -5.123974E-8
+ ppdiblc1 = -5.303252E-14 pdiblc2 = 2.56628E-2 lpdiblc2 = -2.055259E-8
+ wpdiblc2 = -1.714384E-8 ppdiblc2 = 1.490979E-14 pdiblcb = -0.025
+ drout = -1.664994 ldrout = 1.410698E-6 wdrout = 1.516788E-6
+ pdrout = -1.023385E-12 pscbe1 = 2.408892E8 lpscbe1 = 0.261161
+ wpscbe1 = 27.020939 ppscbe1 = -1.894582E-7 pscbe2 = 1.218829E-8
+ lpscbe2 = 1.711727E-15 wpscbe2 = 1.687156E-15 ppscbe2 = -1.241766E-21
+ pvag = 0 delta = 0.01 fprout = 0
+ pdits = 0 pditsl = 0 pditsd = 0
+ lambda = 0 vtl = 0 lc = 5E-9
+ xn = 3 alpha0 = -5.73873E-5 lalpha0 = 4.070202E-11
+ walpha0 = 4.163146E-11 palpha0 = -2.952711E-17 alpha1 = 6.447868E-10
+ lalpha1 = -3.8639E-16 walpha1 = -3.952134E-16 palpha1 = 2.803051E-22
+ beta0 = -199.718245 lbeta0 = 1.437779E-4 wbeta0 = 1.470611E-4
+ pbeta0 = -1.043031E-10 aigbacc = 0.43 bigbacc = 0.054
+ cigbacc = 0.075 nigbacc = 1 aigbinv = 0.35
+ bigbinv = 0.03 cigbinv = 6E-3 eigbinv = 1.1
+ nigbinv = 3 aigc = 0.43 bigc = 0.054
+ cigc = 0.075 aigsd = 0.43 bigsd = 0.054
+ cigsd = 0.075 dlcig = 0 nigc = 1
+ poxedge = 1 pigcd = 1 ntox = 1
+ toxref = 1.175E-8 agidl = 2.626682E-6 lagidl = -2.442578E-12
+ wagidl = -1.905785E-12 pagidl = 1.772273E-18 bgidl = -6.860172E8
+ lbgidl = 734.799841 wbgidl = 1.24379E3 pbgidl = -5.330576E-4
+ cgidl = 2.116464E4 lcgidl = -1.83466E-2 wcgidl = -1.46327E-2
+ pcgidl = 1.330945E-8 egidl = 6.338186 legidl = -4.77685E-6
+ wegidl = -3.938092E-6 pegidl = 3.465347E-12 noia = 3E40
+ noib = 8.53E24 noic = 8.4E7 em = 4.1E7
+ af = 1 ef = 0.88 kf = 0
+ lintnoi = 0 tnoia = 1.5 tnoib = 3.5
+ ntnoi = 1 rnoia = 0.577 rnoib = 0.37
+ xpart = 0 cgso = {1.94171E-10/sw_func_tox_hv_ratio} cgdo = {1.94171E-10/sw_func_tox_hv_ratio}
+ cgbo = {0/sw_func_tox_hv_ratio} ckappas = 0.6 cf = 1.2E-11
+ clc = 1E-7 cle = 0.6 dlc = 4.4983E-8
+ dwc = 0 vfbcv = -0.144689 noff = 4
+ voffcv = 0 acde = 0.401 moin = 15.773
+ cgsl = {9.82591E-12/sw_func_tox_hv_ratio} cgdl = {9.82591E-12/sw_func_tox_hv_ratio} ijthsrev = 0.1
+ ijthsfwd = 0.1 xjbvs = 1 bvs = 12.69
+ jss = 2.1483E-5 jsws = 4.02E-12 cjs = {sw_psd_nw_cj}
+ mjs = 0.33956 mjsws = 0.24676 cjsws = {9.960545E-11*sw_func_psd_nw_cj}
+ cjswgs = {1.47314E-10*sw_func_psd_nw_cj} mjswgs = 0.81 pbs = 0.6587
+ pbsws = 1 pbswgs = 3 xrcrg1 = 12
+ xrcrg2 = 1 rbpb = 50 rbpd = 50
+ rbps = 50 rbdb = 50 rbsb = 50
+ gbmin = 1E-12 tnom = 30 ute = -1.343412
+ lute = -9.673283E-8 kt1 = -0.56587 lkt1 = -8.339359E-8
+ wkt1 = -6.086743E-8 pkt1 = 6.166712E-14 kt1l = 0
+ kt2 = -0.019032 ua1 = 5.524E-10 ub1 = -4.423733E-18
+ wub1 = 6.041755E-25 uc1 = -1.092E-10 at = 2.098824E5
+ lat = -0.141767 wat = -7.90427E-2 pat = 5.606102E-8
+ prt = 0 njs = 1.3632 xtis = 10
+ tpb = 1.671E-3 tpbsw = 0 tpbswg = 0
+ tcj = 9.6E-4 tcjsw = 3E-5 tcjswg = 0
+ tvoff = 0 tvfbsdoff = 0 saref = 2.81E-6
+ sbref = 2.81E-6 wlod = 0 ku0 = 7E-8
+ kvsat = 0.4 kvth0 = 3.5E-8 tku0 = 0
+ llodku0 = 0 wlodku0 = 1 llodvth = 0
+ wlodvth = 1 lku0 = 0 wku0 = 0
+ pku0 = 0 lkvth0 = 0 wkvth0 = 6.5E-7
+ pkvth0 = 0 stk2 = 0 lodk2 = 1
+ steta0 = 0 lodeta0 = 1

.model phv_model.48 pmos
+ level = 54 lmin = 6E-7 lmax = 8E-7 wmin = 4.2E-7
+ wmax = 7.5E-7 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 1.175E-8
+ toxm = 1.175E-8 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 1E23 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {1.2277E-8+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {4.5375E-8-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = -4.7338E-9 dwb = 0 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = -0.745765 lvth0 = -8.277669E-8
+ wvth0 = -7.648133E-8 pvth0 = 3.157951E-14 k1 = 0.782176
+ lk1 = -1.286445E-7 wk1 = -1.103109E-7 pk1 = 5.716581E-14
+ k2 = -8.01078E-2 lk2 = 7.884113E-8 wk2 = 4.938534E-8
+ pk2 = -3.147653E-14 k3 = -2.2405 k3b = -0.172
+ w0 = 0 lpe0 = 0 lpeb = 0
+ vbm = -3 dvtp0 = 0 dvtp1 = 0
+ dvt0 = 4.657 dvt1 = 0.34864 dvt2 = -0.030206
+ dvt0w = -2.2 dvt1w = 1.0163E6 dvt2w = 0
+ vfbsdoff = 0 u0 = 1.32985E-2 lu0 = 9.810583E-10
+ wu0 = 3.244395E-9 pu0 = -1.325881E-15 ua = 2.289509E-9
+ lua = 2.157613E-16 wua = 1.107162E-16 pua = -3.670255E-22
+ ub = -1.772679E-18 lub = 3.613905E-25 wub = 4.960775E-25
+ pub = 1.730732E-31 uc = 1.096683E-11 luc = -8.437516E-18
+ wuc = -5.751589E-18 puc = 3.118473E-24 ud = 0
+ up = 0 lp = 1 eu = 1.67
+ vsat = 5.968524E4 lvsat = 5.805393E-3 wvsat = 6.075244E-4
+ pvsat = 1.935767E-9 a0 = 0.624571 la0 = 5.935088E-8
+ wa0 = 1.883992E-7 pa0 = -1.176269E-13 ags = -2.569696
+ lags = 2.151747E-6 wags = 1.150059E-6 pags = -8.319981E-13
+ b0 = 0 b1 = 0 keta = 8.10983E-2
+ lketa = -8.320234E-8 wketa = -5.444314E-8 pketa = 4.046096E-14
+ a1 = 0 a2 = 0.5 rdsw = 788.47
+ rdswmin = 0 rdw = 0 rdwmin = 0
+ rsw = 0 rswmin = 0 prwb = 0.053538
+ prwg = 0 wr = 1 voff = 9.32315E-2
+ lvoff = -9.065218E-8 wvoff = -7.910169E-8 pvoff = 3.492951E-14
+ voffl = 0 minv = 0 nfactor = 0.265424
+ lnfactor = 1.084101E-6 wnfactor = 8.675217E-7 pnfactor = -6.476487E-13
+ eta0 = -1.894292 leta0 = 9.833736E-7 weta0 = 1.341135E-6
+ peta0 = -6.713485E-13 etab = -0.118866 letab = 7.754305E-8
+ wetab = 8.314016E-8 petab = -5.62947E-14 dsub = -0.142537
+ ldsub = 1.949443E-7 wdsub = 4.181094E-7 pdsub = -2.020606E-13
+ cit = 3.124773E-5 lcit = -1.082041E-11 wcit = -1.541408E-11
+ pcit = 7.849622E-18 cdsc = 0 cdscb = 0
+ cdscd = 0 pclm = 2.438357 lpclm = -7.494714E-7
+ wpclm = -6.765601E-7 ppclm = 3.713441E-13 pdiblc1 = 2.624927
+ lpdiblc1 = -1.35084E-6 wpdiblc1 = -8.31314E-7 ppdiblc1 = 5.002351E-13
+ pdiblc2 = -2.26102E-2 lpdiblc2 = 1.368506E-8 wpdiblc2 = 1.478248E-8
+ ppdiblc2 = -7.733951E-15 pdiblcb = -0.025 drout = -2.257803
+ ldrout = 1.831148E-6 wdrout = 8.862728E-7 pdrout = -5.76192E-13
+ pscbe1 = -2.086815E8 lpscbe1 = 319.119186 wpscbe1 = 128.058083
+ ppscbe1 = -7.185005E-5 pscbe2 = 1.13881E-8 lpscbe2 = 2.279257E-15
+ wpscbe2 = 1.847522E-15 ppscbe2 = -1.355506E-21 pvag = 0
+ delta = 0.01 fprout = 0 pdits = 0
+ pditsl = 0 pditsd = 0 lambda = 0
+ vtl = 0 lc = 5E-9 xn = 3
+ alpha0 = -4.823214E-5 lalpha0 = 3.420872E-11 walpha0 = -9.122915E-13
+ palpha0 = 6.470427E-19 alpha1 = 3.54625E-10 lalpha1 = -1.805928E-16
+ beta0 = -112.746264 lbeta0 = 8.209304E-5 wbeta0 = 3.391603E-6
+ pbeta0 = -2.405495E-12 aigbacc = 0.43 bigbacc = 0.054
+ cigbacc = 0.075 nigbacc = 1 aigbinv = 0.35
+ bigbinv = 0.03 cigbinv = 6E-3 eigbinv = 1.1
+ nigbinv = 3 aigc = 0.43 bigc = 0.054
+ cigc = 0.075 aigsd = 0.43 bigsd = 0.054
+ cigsd = 0.075 dlcig = 0 nigc = 1
+ poxedge = 1 pigcd = 1 ntox = 1
+ toxref = 1.175E-8 agidl = -2.839758E-6 lagidl = 1.434494E-12
+ wagidl = 1.999382E-12 pagidl = -9.974671E-19 bgidl = -3.921719E9
+ lbgidl = 3.029722E3 wbgidl = 2.195213E3 pbgidl = -1.207855E-3
+ cgidl = -1.555729E4 lcgidl = 7.698454E-3 wcgidl = 1.22917E-2
+ pcgidl = -5.786647E-9 egidl = -2.523328 legidl = 1.508179E-6
+ wegidl = 2.454255E-6 pegidl = -1.068426E-12 noia = 3E40
+ noib = 8.53E24 noic = 8.4E7 em = 4.1E7
+ af = 1 ef = 0.88 kf = 0
+ lintnoi = 0 tnoia = 1.5 tnoib = 3.5
+ ntnoi = 1 rnoia = 0.577 rnoib = 0.37
+ xpart = 0 cgso = {1.94171E-10/sw_func_tox_hv_ratio} cgdo = {1.94171E-10/sw_func_tox_hv_ratio}
+ cgbo = {0/sw_func_tox_hv_ratio} ckappas = 0.6 cf = 1.2E-11
+ clc = 1E-7 cle = 0.6 dlc = 4.4983E-8
+ dwc = 0 vfbcv = -0.144689 noff = 4
+ voffcv = 0 acde = 0.401 moin = 15.773
+ cgsl = {9.82591E-12/sw_func_tox_hv_ratio} cgdl = {9.82591E-12/sw_func_tox_hv_ratio} ijthsrev = 0.1
+ ijthsfwd = 0.1 xjbvs = 1 bvs = 12.69
+ jss = 2.1483E-5 jsws = 4.02E-12 cjs = {sw_psd_nw_cj}
+ mjs = 0.33956 mjsws = 0.24676 cjsws = {9.960545E-11*sw_func_psd_nw_cj}
+ cjswgs = {1.47314E-10*sw_func_psd_nw_cj} mjswgs = 0.81 pbs = 0.6587
+ pbsws = 1 pbswgs = 3 xrcrg1 = 12
+ xrcrg2 = 1 rbpb = 50 rbpd = 50
+ rbps = 50 rbdb = 50 rbsb = 50
+ gbmin = 1E-12 tnom = 30 ute = -1.368619
+ lute = -7.885483E-8 wute = -2.842133E-7 pute = 2.015783E-13
+ kt1 = -0.635186 lkt1 = -3.423103E-8 wkt1 = -7.122969E-9
+ pkt1 = 2.354887E-14 kt1l = 0 kt2 = -0.019032
+ ua1 = 5.524E-10 ub1 = -6.399957E-18 lub1 = 1.401637E-24
+ wub1 = 3.522793E-25 pub1 = 1.786574E-31 uc1 = -1.092E-10
+ at = 3.798738E4 lat = -0.01985 wat = -1.10675E-2
+ pat = 7.849622E-9 prt = 0 njs = 1.3632
+ xtis = 10 tpb = 1.671E-3 tpbsw = 0
+ tpbswg = 0 tcj = 9.6E-4 tcjsw = 3E-5
+ tcjswg = 0 tvoff = 0 tvfbsdoff = 0
+ saref = 2.41E-6 sbref = 2.41E-6 wlod = 0
+ ku0 = 7E-8 kvsat = 0.4 kvth0 = 3.5E-8
+ tku0 = 0 llodku0 = 0 wlodku0 = 1
+ llodvth = 0 wlodvth = 1 lku0 = 0
+ wku0 = 0 pku0 = 0 lkvth0 = 0
+ wkvth0 = 6.5E-7 pkvth0 = 0 stk2 = 0
+ lodk2 = 1 steta0 = 0 lodeta0 = 1

.model phv_model.49 pmos
+ level = 54 lmin = 5E-7 lmax = 6E-7 wmin = 4.2E-7
+ wmax = 7.5E-7 version = 4.5
+ binunit = 2 mobmod = 0 capmod = 2
+ rdsmod = 0 igcmod = 0 igbmod = 0
+ rbodymod = 1 trnqsmod = 0 acnqsmod = 0
+ fnoimod = 1 tnoimod = 1 diomod = 1
+ tempmod = 0 permod = 1 geomod = 0
+ rgatemod = 0 epsrox = 3.9 toxe = 1.175E-8
+ toxm = 1.175E-8 dtox = 0 xj = 1.5E-7
+ ndep = 1.7E17 ngate = 1E23 nsd = 1E20
+ rsh = {swx_nrds} rshg = 0.1 phin = 0
+ wint = {1.2277E-8+sw_activecd} wl = 0 wln = 1
+ ww = 0 wwn = 1 wwl = 0
+ lint = {4.5375E-8-sw_polycd} ll = 0 lln = 1
+ lw = 0 lwn = 1 lwl = 0
+ llc = 0 lwc = 0 lwlc = 0
+ wlc = 0 wwc = 0 wwlc = 0
+ dwg = -4.7338E-9 dwb = 0 xl = 0
+ xw = 0 dmcg = 0 dmdg = 0
+ dmcgt = 0 xgw = 0 xgl = 0
+ ngcon = 1 vth0 = -0.730006 lvth0 = -9.080196E-8
+ wvth0 = -1.438204E-7 pvth0 = 6.587192E-14 k1 = 0.382063
+ lk1 = 7.511312E-8 wk1 = 1.089455E-7 pk1 = -5.449051E-14
+ k2 = 0.155805 lk2 = -4.129736E-8 wk2 = -7.125391E-8
+ pk2 = 2.995901E-14 k3 = -2.2405 k3b = -0.172
+ w0 = 0 lpe0 = 0 lpeb = 0
+ vbm = -3 dvtp0 = 0 dvtp1 = 0
+ dvt0 = 4.657 dvt1 = 0.34864 dvt2 = -0.030206
+ dvt0w = -2.2 dvt1w = 1.0163E6 dvt2w = 0
+ vfbsdoff = 0 u0 = 1.49277E-2 lu0 = 1.514166E-10
+ wu0 = 8.564977E-10 pu0 = -1.098445E-16 ua = 9.303429E-9
+ lua = -3.356077E-15 wua = -5.390861E-15 pua = 2.434653E-21
+ ub = -1.414494E-17 lub = 6.661967E-24 wub = 1.032616E-23
+ pub = -4.832897E-30 uc = -1.730147E-11 luc = 5.958116E-18
+ wuc = 8.859631E-18 puc = -4.322291E-24 ud = 0
+ up = 0 lp = 1 eu = 1.67
+ vsat = 9.845805E4 lvsat = -1.39397E-2 wvsat = -1.54488E-2
+ pvsat = 1.011247E-8 a0 = -2.250398 la0 = 1.523429E-6
+ wa0 = 2.127601E-6 pa0 = -1.105166E-12 ags = -0.347211
+ lags = 1.019947E-6 wags = 9.692404E-7 pags = -7.399163E-13
+ b0 = 0 b1 = 0 keta = -0.031617
+ lketa = -2.580207E-8 wketa = -1.174712E-8 pketa = 1.871801E-14
+ a1 = 0 a2 = 0.5 rdsw = 788.47
+ rdswmin = 0 rdw = 0 rdwmin = 0
+ rsw = 0 rswmin = 0 prwb = 0.053538
+ prwg = 0 wr = 1 voff = 6.16317E-2
+ lvoff = -7.455999E-8 wvoff = -1.167251E-7 pvoff = 5.408925E-14
+ voffl = 0 minv = 0 nfactor = 5.766743
+ lnfactor = -1.717446E-6 wnfactor = -2.850815E-6 pnfactor = 1.245914E-12
+ eta0 = -0.405539 leta0 = 2.252265E-7 weta0 = 3.436702E-7
+ peta0 = -1.633897E-13 etab = 0.104773 letab = -3.634525E-8
+ wetab = -7.917936E-8 petab = 2.636652E-14 dsub = 0.170214
+ ldsub = 3.567573E-8 wdsub = 7.215013E-8 pdsub = -2.588082E-14
+ cit = 1E-5 cdsc = 0 cdscb = 0
+ cdscd = 0 pclm = 0.92961 lpclm = 1.885783E-8
+ wpclm = 7.950164E-8 ppclm = -1.368034E-14 pdiblc1 = 0.141036
+ lpdiblc1 = -8.591847E-8 wpdiblc1 = 2.858965E-8 ppdiblc1 = 6.232921E-14
+ pdiblc2 = 0.022596 lpdiblc2 = -9.336207E-9 wpdiblc2 = -1.370424E-8
+ ppdiblc2 = 6.772914E-15 pdiblcb = -0.025 drout = 1.870576
+ ldrout = -2.712292E-7 wdrout = -6.315557E-7 pdrout = 1.967622E-13
+ pscbe1 = 3.066011E8 lpscbe1 = 56.711495 wpscbe1 = 67.755824
+ ppscbe1 = -4.114113E-5 pscbe2 = 2.025541E-8 lpscbe2 = -2.236419E-15
+ wpscbe2 = -4.00011E-15 ppscbe2 = 1.622401E-21 pvag = 0
+ delta = 0.01 fprout = 0 pdits = 0
+ pditsl = 0 pditsd = 0 lambda = 0
+ vtl = 0 lc = 5E-9 xn = 3
+ alpha0 = -2.45509E-5 lalpha0 = 2.214905E-11 walpha0 = 3.191045E-11
+ palpha0 = -1.606794E-17 alpha1 = 0 beta0 = 40.313572
+ lbeta0 = 4.147316E-6 wbeta0 = 4.576011E-6 pbeta0 = -3.008654E-12
+ aigbacc = 0.43 bigbacc = 0.054 cigbacc = 0.075
+ nigbacc = 1 aigbinv = 0.35 bigbinv = 0.03
+ cigbinv = 6E-3 eigbinv = 1.1 nigbinv = 3
+ aigc = 0.43 bigc = 0.054 cigc = 0.075
+ aigsd = 0.43 bigsd = 0.054 cigsd = 0.075
+ dlcig = 0 nigc = 1 poxedge = 1
+ pigcd = 1 ntox = 1 toxref = 1.175E-8
+ agidl = -2.119847E-7 lagidl = 9.630082E-14 wagidl = 1.778682E-13
+ pagidl = -6.986105E-20 bgidl = 2.468875E9 lbgidl = -224.688351
+ wbgidl = -496.69448 pbgidl = 1.629993E-4 cgidl = -6.03198E3
+ lcgidl = 2.847692E-3 wcgidl = 4.985251E-3 pcgidl = -2.065847E-9
+ egidl = -0.475833 legidl = 4.654919E-7 wegidl = 1.019329E-6
+ pegidl = -3.376892E-13 noia = 3E40 noib = 8.53E24
+ noic = 8.4E7 em = 4.1E7 af = 1
+ ef = 0.88 kf = 0 lintnoi = 0
+ tnoia = 1.5 tnoib = 3.5 ntnoi = 1
+ rnoia = 0.577 rnoib = 0.37 xpart = 0
+ cgso = {1.94171E-10/sw_func_tox_hv_ratio} cgdo = {1.94171E-10/sw_func_tox_hv_ratio} cgbo = {0/sw_func_tox_hv_ratio}
+ ckappas = 0.6 cf = 1.2E-11 clc = 1E-7
+ cle = 0.6 dlc = 4.4983E-8 dwc = 0
+ vfbcv = -0.144689 noff = 4 voffcv = 0
+ acde = 0.401 moin = 15.773 cgsl = {9.82591E-12/sw_func_tox_hv_ratio}
+ cgdl = {9.82591E-12/sw_func_tox_hv_ratio} ijthsrev = 0.1 ijthsfwd = 0.1
+ xjbvs = 1 bvs = 12.69 jss = 2.1483E-5
+ jsws = 4.02E-12 cjs = {sw_psd_nw_cj} mjs = 0.33956
+ mjsws = 0.24676 cjsws = {9.960545E-11*sw_func_psd_nw_cj} cjswgs = {1.47314E-10*sw_func_psd_nw_cj}
+ mjswgs = 0.81 pbs = 0.6587 pbsws = 1
+ pbswgs = 3 xrcrg1 = 12 xrcrg2 = 1
+ rbpb = 50 rbpd = 50 rbps = 50
+ rbdb = 50 rbsb = 50 gbmin = 1E-12
+ tnom = 30 ute = -2.117845 lute = 3.026883E-7
+ wute = 5.428113E-7 pute = -2.19584E-13 kt1 = -0.927994
+ lkt1 = 1.148817E-7 wkt1 = 2.027726E-7 pkt1 = -8.334046E-14
+ kt1l = 0 kt2 = -0.019032 ua1 = 5.52E-10
+ ub1 = -8.671393E-18 lub1 = 2.558365E-24 wub1 = 4.347592E-24
+ pub1 = -1.855956E-30 uc1 = 2.228292E-10 luc1 = -1.690859E-16
+ wuc1 = -2.408692E-16 puc1 = 1.226627E-22 at = 3.824143E4
+ lat = -1.99794E-2 wat = -2.41149E-2 pat = 1.449399E-8
+ prt = 0 njs = 1.3632 xtis = 10
+ tpb = 1.671E-3 tpbsw = 0 tpbswg = 0
+ tcj = 9.6E-4 tcjsw = 3E-5 tcjswg = 0
+ tvoff = 0 tvfbsdoff = 0 saref = 2.02E-6
+ sbref = 2.01E-6 wlod = 0 ku0 = 7E-8
+ kvsat = 0.4 kvth0 = 3.5E-8 tku0 = 0
+ llodku0 = 0 wlodku0 = 1 llodvth = 0
+ wlodvth = 1 lku0 = 0 wku0 = 0
+ pku0 = 0 lkvth0 = 0 wkvth0 = 6.5E-7
+ pkvth0 = 0 stk2 = 0 lodk2 = 1
+ steta0 = 0 lodeta0 = 1

.ends sky130_fd_pr__pfet_g5v0d10v5
